netcdf test_proleptic_gregorian {
dimensions:
	time = UNLIMITED ;
	lat = 2 ;
	lon = 2 ;
    bnds = 2 ;
variables:
	double time(time) ;
		time:bounds = "time_bnds" ;
		time:units = "days since 0001-01-01" ;
		time:calendar = "proleptic_gregorian" ;
		time:axis = "T" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
	double time_bnds(time, bnds) ;
	float lat ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "Latitude" ;
	float lon ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "Longitude" ;
	float z ;
		z:standard_name = "depth" ;
		z:positive = "down" ;
		z:units = "m" ;
		z:long_name = "Depth below surface" ;
	float temperature(time, lat, lon) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "deg_C" ;
		temperature:long_name = "Seawater Temperature" ;
		temperature:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:variable_id = "temp-max" ;
		:scenario = "sres-a1b" ;
		:dataset_id = "ukcp18-land-prob-25km" ;
		:prob_type = "sample" ;
		:frequency = "mon" ;
data:

 time = 675348.5, 675378, 675407.5, 675438, 675468.5, 675499, 675529.5,
    675560.5, 675591, 675621.5, 675652, 675682.5, 675713.5, 675743, 675772.5,
    675803, 675833.5, 675864, 675894.5, 675925.5, 675956, 675986.5, 676017,
    676047.5, 676078.5, 676108.5, 676138.5, 676169, 676199.5, 676230,
    676260.5, 676291.5, 676322, 676352.5, 676383, 676413.5, 676444.5, 676474,
    676503.5, 676534, 676564.5, 676595, 676625.5, 676656.5, 676687, 676717.5,
    676748, 676778.5, 676809.5, 676839, 676868.5, 676899, 676929.5, 676960,
    676990.5, 677021.5, 677052, 677082.5, 677113, 677143.5, 677174.5, 677204,
    677233.5, 677264, 677294.5, 677325, 677355.5, 677386.5, 677417, 677447.5,
    677478, 677508.5, 677539.5, 677569.5, 677599.5, 677630, 677660.5, 677691,
    677721.5, 677752.5, 677783, 677813.5, 677844, 677874.5, 677905.5, 677935,
    677964.5, 677995, 678025.5, 678056, 678086.5, 678117.5, 678148, 678178.5,
    678209, 678239.5, 678270.5, 678300, 678329.5, 678360, 678390.5, 678421,
    678451.5, 678482.5, 678513, 678543.5, 678574, 678604.5, 678635.5, 678665,
    678694.5, 678725, 678755.5, 678786, 678816.5, 678847.5, 678878, 678908.5,
    678939, 678969.5, 679000.5, 679030.5, 679060.5, 679091, 679121.5, 679152,
    679182.5, 679213.5, 679244, 679274.5, 679305, 679335.5, 679366.5, 679396,
    679425.5, 679456, 679486.5, 679517, 679547.5, 679578.5, 679609, 679639.5,
    679670, 679700.5, 679731.5, 679761, 679790.5, 679821, 679851.5, 679882,
    679912.5, 679943.5, 679974, 680004.5, 680035, 680065.5, 680096.5, 680126,
    680155.5, 680186, 680216.5, 680247, 680277.5, 680308.5, 680339, 680369.5,
    680400, 680430.5, 680461.5, 680491.5, 680521.5, 680552, 680582.5, 680613,
    680643.5, 680674.5, 680705, 680735.5, 680766, 680796.5, 680827.5, 680857,
    680886.5, 680917, 680947.5, 680978, 681008.5, 681039.5, 681070, 681100.5,
    681131, 681161.5, 681192.5, 681222, 681251.5, 681282, 681312.5, 681343,
    681373.5, 681404.5, 681435, 681465.5, 681496, 681526.5, 681557.5, 681587,
    681616.5, 681647, 681677.5, 681708, 681738.5, 681769.5, 681800, 681830.5,
    681861, 681891.5, 681922.5, 681952.5, 681982.5, 682013, 682043.5, 682074,
    682104.5, 682135.5, 682166, 682196.5, 682227, 682257.5, 682288.5, 682318,
    682347.5, 682378, 682408.5, 682439, 682469.5, 682500.5, 682531, 682561.5,
    682592, 682622.5, 682653.5, 682683, 682712.5, 682743, 682773.5, 682804,
    682834.5, 682865.5, 682896, 682926.5, 682957, 682987.5, 683018.5, 683048,
    683077.5, 683108, 683138.5, 683169, 683199.5, 683230.5, 683261, 683291.5,
    683322, 683352.5, 683383.5, 683413.5, 683443.5, 683474, 683504.5, 683535,
    683565.5, 683596.5, 683627, 683657.5, 683688, 683718.5, 683749.5, 683779,
    683808.5, 683839, 683869.5, 683900, 683930.5, 683961.5, 683992, 684022.5,
    684053, 684083.5, 684114.5, 684144, 684173.5, 684204, 684234.5, 684265,
    684295.5, 684326.5, 684357, 684387.5, 684418, 684448.5, 684479.5, 684509,
    684538.5, 684569, 684599.5, 684630, 684660.5, 684691.5, 684722, 684752.5,
    684783, 684813.5, 684844.5, 684874.5, 684904.5, 684935, 684965.5, 684996,
    685026.5, 685057.5, 685088, 685118.5, 685149, 685179.5, 685210.5, 685240,
    685269.5, 685300, 685330.5, 685361, 685391.5, 685422.5, 685453, 685483.5,
    685514, 685544.5, 685575.5, 685605, 685634.5, 685665, 685695.5, 685726,
    685756.5, 685787.5, 685818, 685848.5, 685879, 685909.5, 685940.5, 685970,
    685999.5, 686030, 686060.5, 686091, 686121.5, 686152.5, 686183, 686213.5,
    686244, 686274.5, 686305.5, 686335.5, 686365.5, 686396, 686426.5, 686457,
    686487.5, 686518.5, 686549, 686579.5, 686610, 686640.5, 686671.5, 686701,
    686730.5, 686761, 686791.5, 686822, 686852.5, 686883.5, 686914, 686944.5,
    686975, 687005.5, 687036.5, 687066, 687095.5, 687126, 687156.5, 687187,
    687217.5, 687248.5, 687279, 687309.5, 687340, 687370.5, 687401.5, 687431,
    687460.5, 687491, 687521.5, 687552, 687582.5, 687613.5, 687644, 687674.5,
    687705, 687735.5, 687766.5, 687796.5, 687826.5, 687857, 687887.5, 687918,
    687948.5, 687979.5, 688010, 688040.5, 688071, 688101.5, 688132.5, 688162,
    688191.5, 688222, 688252.5, 688283, 688313.5, 688344.5, 688375, 688405.5,
    688436, 688466.5, 688497.5, 688527, 688556.5, 688587, 688617.5, 688648,
    688678.5, 688709.5, 688740, 688770.5, 688801, 688831.5, 688862.5, 688892,
    688921.5, 688952, 688982.5, 689013, 689043.5, 689074.5, 689105, 689135.5,
    689166, 689196.5, 689227.5, 689257.5, 689287.5, 689318, 689348.5, 689379,
    689409.5, 689440.5, 689471, 689501.5, 689532, 689562.5, 689593.5, 689623,
    689652.5, 689683, 689713.5, 689744, 689774.5, 689805.5, 689836, 689866.5,
    689897, 689927.5, 689958.5, 689988, 690017.5, 690048, 690078.5, 690109,
    690139.5, 690170.5, 690201, 690231.5, 690262, 690292.5, 690323.5, 690353,
    690382.5, 690413, 690443.5, 690474, 690504.5, 690535.5, 690566, 690596.5,
    690627, 690657.5, 690688.5, 690718.5, 690748.5, 690779, 690809.5, 690840,
    690870.5, 690901.5, 690932, 690962.5, 690993, 691023.5, 691054.5, 691084,
    691113.5, 691144, 691174.5, 691205, 691235.5, 691266.5, 691297, 691327.5,
    691358, 691388.5, 691419.5, 691449, 691478.5, 691509, 691539.5, 691570,
    691600.5, 691631.5, 691662, 691692.5, 691723, 691753.5, 691784.5, 691814,
    691843.5, 691874, 691904.5, 691935, 691965.5, 691996.5, 692027, 692057.5,
    692088, 692118.5, 692149.5, 692179.5, 692209.5, 692240, 692270.5, 692301,
    692331.5, 692362.5, 692393, 692423.5, 692454, 692484.5, 692515.5, 692545,
    692574.5, 692605, 692635.5, 692666, 692696.5, 692727.5, 692758, 692788.5,
    692819, 692849.5, 692880.5, 692910, 692939.5, 692970, 693000.5, 693031,
    693061.5, 693092.5, 693123, 693153.5, 693184, 693214.5, 693245.5, 693275,
    693304.5, 693335, 693365.5, 693396, 693426.5, 693457.5, 693488, 693518.5,
    693549, 693579.5, 693610.5, 693640, 693669.5, 693700, 693730.5, 693761,
    693791.5, 693822.5, 693853, 693883.5, 693914, 693944.5, 693975.5, 694005,
    694034.5, 694065, 694095.5, 694126, 694156.5, 694187.5, 694218, 694248.5,
    694279, 694309.5, 694340.5, 694370, 694399.5, 694430, 694460.5, 694491,
    694521.5, 694552.5, 694583, 694613.5, 694644, 694674.5, 694705.5, 694735,
    694764.5, 694795, 694825.5, 694856, 694886.5, 694917.5, 694948, 694978.5,
    695009, 695039.5, 695070.5, 695100.5, 695130.5, 695161, 695191.5, 695222,
    695252.5, 695283.5, 695314, 695344.5, 695375, 695405.5, 695436.5, 695466,
    695495.5, 695526, 695556.5, 695587, 695617.5, 695648.5, 695679, 695709.5,
    695740, 695770.5, 695801.5, 695831, 695860.5, 695891, 695921.5, 695952,
    695982.5, 696013.5, 696044, 696074.5, 696105, 696135.5, 696166.5, 696196,
    696225.5, 696256, 696286.5, 696317, 696347.5, 696378.5, 696409, 696439.5,
    696470, 696500.5, 696531.5, 696561.5, 696591.5, 696622, 696652.5, 696683,
    696713.5, 696744.5, 696775, 696805.5, 696836, 696866.5, 696897.5, 696927,
    696956.5, 696987, 697017.5, 697048, 697078.5, 697109.5, 697140, 697170.5,
    697201, 697231.5, 697262.5, 697292, 697321.5, 697352, 697382.5, 697413,
    697443.5, 697474.5, 697505, 697535.5, 697566, 697596.5, 697627.5, 697657,
    697686.5, 697717, 697747.5, 697778, 697808.5, 697839.5, 697870, 697900.5,
    697931, 697961.5, 697992.5, 698022.5, 698052.5, 698083, 698113.5, 698144,
    698174.5, 698205.5, 698236, 698266.5, 698297, 698327.5, 698358.5, 698388,
    698417.5, 698448, 698478.5, 698509, 698539.5, 698570.5, 698601, 698631.5,
    698662, 698692.5, 698723.5, 698753, 698782.5, 698813, 698843.5, 698874,
    698904.5, 698935.5, 698966, 698996.5, 699027, 699057.5, 699088.5, 699118,
    699147.5, 699178, 699208.5, 699239, 699269.5, 699300.5, 699331, 699361.5,
    699392, 699422.5, 699453.5, 699483.5, 699513.5, 699544, 699574.5, 699605,
    699635.5, 699666.5, 699697, 699727.5, 699758, 699788.5, 699819.5, 699849,
    699878.5, 699909, 699939.5, 699970, 700000.5, 700031.5, 700062, 700092.5,
    700123, 700153.5, 700184.5, 700214, 700243.5, 700274, 700304.5, 700335,
    700365.5, 700396.5, 700427, 700457.5, 700488, 700518.5, 700549.5, 700579,
    700608.5, 700639, 700669.5, 700700, 700730.5, 700761.5, 700792, 700822.5,
    700853, 700883.5, 700914.5, 700944.5, 700974.5, 701005, 701035.5, 701066,
    701096.5, 701127.5, 701158, 701188.5, 701219, 701249.5, 701280.5, 701310,
    701339.5, 701370, 701400.5, 701431, 701461.5, 701492.5, 701523, 701553.5,
    701584, 701614.5, 701645.5, 701675, 701704.5, 701735, 701765.5, 701796,
    701826.5, 701857.5, 701888, 701918.5, 701949, 701979.5, 702010.5, 702040,
    702069.5, 702100, 702130.5, 702161, 702191.5, 702222.5, 702253, 702283.5,
    702314, 702344.5, 702375.5, 702405.5, 702435.5, 702466, 702496.5, 702527,
    702557.5, 702588.5, 702619, 702649.5, 702680, 702710.5, 702741.5, 702771,
    702800.5, 702831, 702861.5, 702892, 702922.5, 702953.5, 702984, 703014.5,
    703045, 703075.5, 703106.5, 703136, 703165.5, 703196, 703226.5, 703257,
    703287.5, 703318.5, 703349, 703379.5, 703410, 703440.5, 703471.5, 703501,
    703530.5, 703561, 703591.5, 703622, 703652.5, 703683.5, 703714, 703744.5,
    703775, 703805.5, 703836.5, 703866.5, 703896.5, 703927, 703957.5, 703988,
    704018.5, 704049.5, 704080, 704110.5, 704141, 704171.5, 704202.5, 704232,
    704261.5, 704292, 704322.5, 704353, 704383.5, 704414.5, 704445, 704475.5,
    704506, 704536.5, 704567.5, 704597, 704626.5, 704657, 704687.5, 704718,
    704748.5, 704779.5, 704810, 704840.5, 704871, 704901.5, 704932.5, 704962,
    704991.5, 705022, 705052.5, 705083, 705113.5, 705144.5, 705175, 705205.5,
    705236, 705266.5, 705297.5, 705327.5, 705357.5, 705388, 705418.5, 705449,
    705479.5, 705510.5, 705541, 705571.5, 705602, 705632.5, 705663.5, 705693,
    705722.5, 705753, 705783.5, 705814, 705844.5, 705875.5, 705906, 705936.5,
    705967, 705997.5, 706028.5, 706058, 706087.5, 706118, 706148.5, 706179,
    706209.5, 706240.5, 706271, 706301.5, 706332, 706362.5, 706393.5, 706423,
    706452.5, 706483, 706513.5, 706544, 706574.5, 706605.5, 706636, 706666.5,
    706697, 706727.5, 706758.5, 706788.5, 706818.5, 706849, 706879.5, 706910,
    706940.5, 706971.5, 707002, 707032.5, 707063, 707093.5, 707124.5, 707154,
    707183.5, 707214, 707244.5, 707275, 707305.5, 707336.5, 707367, 707397.5,
    707428, 707458.5, 707489.5, 707519, 707548.5, 707579, 707609.5, 707640,
    707670.5, 707701.5, 707732, 707762.5, 707793, 707823.5, 707854.5, 707884,
    707913.5, 707944, 707974.5, 708005, 708035.5, 708066.5, 708097, 708127.5,
    708158, 708188.5, 708219.5, 708249.5, 708279.5, 708310, 708340.5, 708371,
    708401.5, 708432.5, 708463, 708493.5, 708524, 708554.5, 708585.5, 708615,
    708644.5, 708675, 708705.5, 708736, 708766.5, 708797.5, 708828, 708858.5,
    708889, 708919.5, 708950.5, 708980, 709009.5, 709040, 709070.5, 709101,
    709131.5, 709162.5, 709193, 709223.5, 709254, 709284.5, 709315.5, 709345,
    709374.5, 709405, 709435.5, 709466, 709496.5, 709527.5, 709558, 709588.5,
    709619, 709649.5, 709680.5, 709710.5, 709740.5, 709771, 709801.5, 709832,
    709862.5, 709893.5, 709924, 709954.5, 709985, 710015.5, 710046.5, 710076,
    710105.5, 710136, 710166.5, 710197, 710227.5, 710258.5, 710289, 710319.5,
    710350, 710380.5, 710411.5, 710441, 710470.5, 710501, 710531.5, 710562,
    710592.5, 710623.5, 710654, 710684.5, 710715, 710745.5, 710776.5, 710806,
    710835.5, 710866, 710896.5, 710927, 710957.5, 710988.5, 711019, 711049.5,
    711080, 711110.5, 711141.5, 711171.5, 711201.5, 711232, 711262.5, 711293,
    711323.5, 711354.5, 711385, 711415.5, 711446, 711476.5, 711507.5, 711537,
    711566.5, 711597, 711627.5, 711658, 711688.5, 711719.5, 711750, 711780.5,
    711811, 711841.5, 711872.5, 711902, 711931.5, 711962, 711992.5, 712023,
    712053.5, 712084.5, 712115, 712145.5, 712176, 712206.5, 712237.5, 712267,
    712296.5, 712327, 712357.5, 712388, 712418.5, 712449.5, 712480, 712510.5,
    712541, 712571.5, 712602.5, 712632.5, 712662.5, 712693, 712723.5, 712754,
    712784.5, 712815.5, 712846, 712876.5, 712907, 712937.5, 712968.5, 712998,
    713027.5, 713058, 713088.5, 713119, 713149.5, 713180.5, 713211, 713241.5,
    713272, 713302.5, 713333.5, 713363, 713392.5, 713423, 713453.5, 713484,
    713514.5, 713545.5, 713576, 713606.5, 713637, 713667.5, 713698.5, 713728,
    713757.5, 713788, 713818.5, 713849, 713879.5, 713910.5, 713941, 713971.5,
    714002, 714032.5, 714063.5, 714093.5, 714123.5, 714154, 714184.5, 714215,
    714245.5, 714276.5, 714307, 714337.5, 714368, 714398.5, 714429.5, 714459,
    714488.5, 714519, 714549.5, 714580, 714610.5, 714641.5, 714672, 714702.5,
    714733, 714763.5, 714794.5, 714824, 714853.5, 714884, 714914.5, 714945,
    714975.5, 715006.5, 715037, 715067.5, 715098, 715128.5, 715159.5, 715189,
    715218.5, 715249, 715279.5, 715310, 715340.5, 715371.5, 715402, 715432.5,
    715463, 715493.5, 715524.5, 715554.5, 715584.5, 715615, 715645.5, 715676,
    715706.5, 715737.5, 715768, 715798.5, 715829, 715859.5, 715890.5, 715920,
    715949.5, 715980, 716010.5, 716041, 716071.5, 716102.5, 716133, 716163.5,
    716194, 716224.5, 716255.5, 716285, 716314.5, 716345, 716375.5, 716406,
    716436.5, 716467.5, 716498, 716528.5, 716559, 716589.5, 716620.5, 716650,
    716679.5, 716710, 716740.5, 716771, 716801.5, 716832.5, 716863, 716893.5,
    716924, 716954.5, 716985.5, 717015.5, 717045.5, 717076, 717106.5, 717137,
    717167.5, 717198.5, 717229, 717259.5, 717290, 717320.5, 717351.5, 717381,
    717410.5, 717441, 717471.5, 717502, 717532.5, 717563.5, 717594, 717624.5,
    717655, 717685.5, 717716.5, 717746, 717775.5, 717806, 717836.5, 717867,
    717897.5, 717928.5, 717959, 717989.5, 718020, 718050.5, 718081.5, 718111,
    718140.5, 718171, 718201.5, 718232, 718262.5, 718293.5, 718324, 718354.5,
    718385, 718415.5, 718446.5, 718476.5, 718506.5, 718537, 718567.5, 718598,
    718628.5, 718659.5, 718690, 718720.5, 718751, 718781.5, 718812.5, 718842,
    718871.5, 718902, 718932.5, 718963, 718993.5, 719024.5, 719055, 719085.5,
    719116, 719146.5, 719177.5, 719207, 719236.5, 719267, 719297.5, 719328,
    719358.5, 719389.5, 719420, 719450.5, 719481, 719511.5, 719542.5, 719572,
    719601.5, 719632, 719662.5, 719693, 719723.5, 719754.5, 719785, 719815.5,
    719846, 719876.5, 719907.5, 719937.5, 719967.5, 719998, 720028.5, 720059,
    720089.5, 720120.5, 720151, 720181.5, 720212, 720242.5, 720273.5, 720303,
    720332.5, 720363, 720393.5, 720424, 720454.5, 720485.5, 720516, 720546.5,
    720577, 720607.5, 720638.5, 720668, 720697.5, 720728, 720758.5, 720789,
    720819.5, 720850.5, 720881, 720911.5, 720942, 720972.5, 721003.5, 721033,
    721062.5, 721093, 721123.5, 721154, 721184.5, 721215.5, 721246, 721276.5,
    721307, 721337.5, 721368.5, 721398.5, 721428.5, 721459, 721489.5, 721520,
    721550.5, 721581.5, 721612, 721642.5, 721673, 721703.5, 721734.5, 721764,
    721793.5, 721824, 721854.5, 721885, 721915.5, 721946.5, 721977, 722007.5,
    722038, 722068.5, 722099.5, 722129, 722158.5, 722189, 722219.5, 722250,
    722280.5, 722311.5, 722342, 722372.5, 722403, 722433.5, 722464.5, 722494,
    722523.5, 722554, 722584.5, 722615, 722645.5, 722676.5, 722707, 722737.5,
    722768, 722798.5, 722829.5, 722859.5, 722889.5, 722920, 722950.5, 722981,
    723011.5, 723042.5, 723073, 723103.5, 723134, 723164.5, 723195.5, 723225,
    723254.5, 723285, 723315.5, 723346, 723376.5, 723407.5, 723438, 723468.5,
    723499, 723529.5, 723560.5, 723590, 723619.5, 723650, 723680.5, 723711,
    723741.5, 723772.5, 723803, 723833.5, 723864, 723894.5, 723925.5, 723955,
    723984.5, 724015, 724045.5, 724076, 724106.5, 724137.5, 724168, 724198.5,
    724229, 724259.5, 724290.5, 724320.5, 724350.5, 724381, 724411.5, 724442,
    724472.5, 724503.5, 724534, 724564.5, 724595, 724625.5, 724656.5, 724686,
    724715.5, 724746, 724776.5, 724807, 724837.5, 724868.5, 724899, 724929.5,
    724960, 724990.5, 725021.5, 725051, 725080.5, 725111, 725141.5, 725172,
    725202.5, 725233.5, 725264, 725294.5, 725325, 725355.5, 725386.5, 725416,
    725445.5, 725476, 725506.5, 725537, 725567.5, 725598.5, 725629, 725659.5,
    725690, 725720.5, 725751.5, 725781.5, 725811.5, 725842, 725872.5, 725903,
    725933.5, 725964.5, 725995, 726025.5, 726056, 726086.5, 726117.5, 726147,
    726176.5, 726207, 726237.5, 726268, 726298.5, 726329.5, 726360, 726390.5,
    726421, 726451.5, 726482.5, 726512, 726541.5, 726572, 726602.5, 726633,
    726663.5, 726694.5, 726725, 726755.5, 726786, 726816.5, 726847.5, 726877,
    726906.5, 726937, 726967.5, 726998, 727028.5, 727059.5, 727090, 727120.5,
    727151, 727181.5, 727212.5, 727242.5, 727272.5, 727303, 727333.5, 727364,
    727394.5, 727425.5, 727456, 727486.5, 727517, 727547.5, 727578.5, 727608,
    727637.5, 727668, 727698.5, 727729, 727759.5, 727790.5, 727821, 727851.5,
    727882, 727912.5, 727943.5, 727973, 728002.5, 728033, 728063.5, 728094,
    728124.5, 728155.5, 728186, 728216.5, 728247, 728277.5, 728308.5, 728338,
    728367.5, 728398, 728428.5, 728459, 728489.5, 728520.5, 728551, 728581.5,
    728612, 728642.5, 728673.5, 728703.5, 728733.5, 728764, 728794.5, 728825,
    728855.5, 728886.5, 728917, 728947.5, 728978, 729008.5, 729039.5, 729069,
    729098.5, 729129, 729159.5, 729190, 729220.5, 729251.5, 729282, 729312.5,
    729343, 729373.5, 729404.5, 729434, 729463.5, 729494, 729524.5, 729555,
    729585.5, 729616.5, 729647, 729677.5, 729708, 729738.5, 729769.5, 729799,
    729828.5, 729859, 729889.5, 729920, 729950.5, 729981.5, 730012, 730042.5,
    730073, 730103.5, 730134.5, 730164.5, 730194.5, 730225, 730255.5, 730286,
    730316.5, 730347.5, 730378, 730408.5, 730439, 730469.5, 730500.5, 730530,
    730559.5, 730590, 730620.5, 730651, 730681.5, 730712.5, 730743, 730773.5,
    730804, 730834.5, 730865.5, 730895, 730924.5, 730955, 730985.5, 731016,
    731046.5, 731077.5, 731108, 731138.5, 731169, 731199.5, 731230.5, 731260,
    731289.5, 731320, 731350.5, 731381, 731411.5, 731442.5, 731473, 731503.5,
    731534, 731564.5, 731595.5, 731625.5, 731655.5, 731686, 731716.5, 731747,
    731777.5, 731808.5, 731839, 731869.5, 731900, 731930.5, 731961.5, 731991,
    732020.5, 732051, 732081.5, 732112, 732142.5, 732173.5, 732204, 732234.5,
    732265, 732295.5 ;

 time_bnds =
  675333, 675364,
  675364, 675392,
  675392, 675423,
  675423, 675453,
  675453, 675484,
  675484, 675514,
  675514, 675545,
  675545, 675576,
  675576, 675606,
  675606, 675637,
  675637, 675667,
  675667, 675698,
  675698, 675729,
  675729, 675757,
  675757, 675788,
  675788, 675818,
  675818, 675849,
  675849, 675879,
  675879, 675910,
  675910, 675941,
  675941, 675971,
  675971, 676002,
  676002, 676032,
  676032, 676063,
  676063, 676094,
  676094, 676123,
  676123, 676154,
  676154, 676184,
  676184, 676215,
  676215, 676245,
  676245, 676276,
  676276, 676307,
  676307, 676337,
  676337, 676368,
  676368, 676398,
  676398, 676429,
  676429, 676460,
  676460, 676488,
  676488, 676519,
  676519, 676549,
  676549, 676580,
  676580, 676610,
  676610, 676641,
  676641, 676672,
  676672, 676702,
  676702, 676733,
  676733, 676763,
  676763, 676794,
  676794, 676825,
  676825, 676853,
  676853, 676884,
  676884, 676914,
  676914, 676945,
  676945, 676975,
  676975, 677006,
  677006, 677037,
  677037, 677067,
  677067, 677098,
  677098, 677128,
  677128, 677159,
  677159, 677190,
  677190, 677218,
  677218, 677249,
  677249, 677279,
  677279, 677310,
  677310, 677340,
  677340, 677371,
  677371, 677402,
  677402, 677432,
  677432, 677463,
  677463, 677493,
  677493, 677524,
  677524, 677555,
  677555, 677584,
  677584, 677615,
  677615, 677645,
  677645, 677676,
  677676, 677706,
  677706, 677737,
  677737, 677768,
  677768, 677798,
  677798, 677829,
  677829, 677859,
  677859, 677890,
  677890, 677921,
  677921, 677949,
  677949, 677980,
  677980, 678010,
  678010, 678041,
  678041, 678071,
  678071, 678102,
  678102, 678133,
  678133, 678163,
  678163, 678194,
  678194, 678224,
  678224, 678255,
  678255, 678286,
  678286, 678314,
  678314, 678345,
  678345, 678375,
  678375, 678406,
  678406, 678436,
  678436, 678467,
  678467, 678498,
  678498, 678528,
  678528, 678559,
  678559, 678589,
  678589, 678620,
  678620, 678651,
  678651, 678679,
  678679, 678710,
  678710, 678740,
  678740, 678771,
  678771, 678801,
  678801, 678832,
  678832, 678863,
  678863, 678893,
  678893, 678924,
  678924, 678954,
  678954, 678985,
  678985, 679016,
  679016, 679045,
  679045, 679076,
  679076, 679106,
  679106, 679137,
  679137, 679167,
  679167, 679198,
  679198, 679229,
  679229, 679259,
  679259, 679290,
  679290, 679320,
  679320, 679351,
  679351, 679382,
  679382, 679410,
  679410, 679441,
  679441, 679471,
  679471, 679502,
  679502, 679532,
  679532, 679563,
  679563, 679594,
  679594, 679624,
  679624, 679655,
  679655, 679685,
  679685, 679716,
  679716, 679747,
  679747, 679775,
  679775, 679806,
  679806, 679836,
  679836, 679867,
  679867, 679897,
  679897, 679928,
  679928, 679959,
  679959, 679989,
  679989, 680020,
  680020, 680050,
  680050, 680081,
  680081, 680112,
  680112, 680140,
  680140, 680171,
  680171, 680201,
  680201, 680232,
  680232, 680262,
  680262, 680293,
  680293, 680324,
  680324, 680354,
  680354, 680385,
  680385, 680415,
  680415, 680446,
  680446, 680477,
  680477, 680506,
  680506, 680537,
  680537, 680567,
  680567, 680598,
  680598, 680628,
  680628, 680659,
  680659, 680690,
  680690, 680720,
  680720, 680751,
  680751, 680781,
  680781, 680812,
  680812, 680843,
  680843, 680871,
  680871, 680902,
  680902, 680932,
  680932, 680963,
  680963, 680993,
  680993, 681024,
  681024, 681055,
  681055, 681085,
  681085, 681116,
  681116, 681146,
  681146, 681177,
  681177, 681208,
  681208, 681236,
  681236, 681267,
  681267, 681297,
  681297, 681328,
  681328, 681358,
  681358, 681389,
  681389, 681420,
  681420, 681450,
  681450, 681481,
  681481, 681511,
  681511, 681542,
  681542, 681573,
  681573, 681601,
  681601, 681632,
  681632, 681662,
  681662, 681693,
  681693, 681723,
  681723, 681754,
  681754, 681785,
  681785, 681815,
  681815, 681846,
  681846, 681876,
  681876, 681907,
  681907, 681938,
  681938, 681967,
  681967, 681998,
  681998, 682028,
  682028, 682059,
  682059, 682089,
  682089, 682120,
  682120, 682151,
  682151, 682181,
  682181, 682212,
  682212, 682242,
  682242, 682273,
  682273, 682304,
  682304, 682332,
  682332, 682363,
  682363, 682393,
  682393, 682424,
  682424, 682454,
  682454, 682485,
  682485, 682516,
  682516, 682546,
  682546, 682577,
  682577, 682607,
  682607, 682638,
  682638, 682669,
  682669, 682697,
  682697, 682728,
  682728, 682758,
  682758, 682789,
  682789, 682819,
  682819, 682850,
  682850, 682881,
  682881, 682911,
  682911, 682942,
  682942, 682972,
  682972, 683003,
  683003, 683034,
  683034, 683062,
  683062, 683093,
  683093, 683123,
  683123, 683154,
  683154, 683184,
  683184, 683215,
  683215, 683246,
  683246, 683276,
  683276, 683307,
  683307, 683337,
  683337, 683368,
  683368, 683399,
  683399, 683428,
  683428, 683459,
  683459, 683489,
  683489, 683520,
  683520, 683550,
  683550, 683581,
  683581, 683612,
  683612, 683642,
  683642, 683673,
  683673, 683703,
  683703, 683734,
  683734, 683765,
  683765, 683793,
  683793, 683824,
  683824, 683854,
  683854, 683885,
  683885, 683915,
  683915, 683946,
  683946, 683977,
  683977, 684007,
  684007, 684038,
  684038, 684068,
  684068, 684099,
  684099, 684130,
  684130, 684158,
  684158, 684189,
  684189, 684219,
  684219, 684250,
  684250, 684280,
  684280, 684311,
  684311, 684342,
  684342, 684372,
  684372, 684403,
  684403, 684433,
  684433, 684464,
  684464, 684495,
  684495, 684523,
  684523, 684554,
  684554, 684584,
  684584, 684615,
  684615, 684645,
  684645, 684676,
  684676, 684707,
  684707, 684737,
  684737, 684768,
  684768, 684798,
  684798, 684829,
  684829, 684860,
  684860, 684889,
  684889, 684920,
  684920, 684950,
  684950, 684981,
  684981, 685011,
  685011, 685042,
  685042, 685073,
  685073, 685103,
  685103, 685134,
  685134, 685164,
  685164, 685195,
  685195, 685226,
  685226, 685254,
  685254, 685285,
  685285, 685315,
  685315, 685346,
  685346, 685376,
  685376, 685407,
  685407, 685438,
  685438, 685468,
  685468, 685499,
  685499, 685529,
  685529, 685560,
  685560, 685591,
  685591, 685619,
  685619, 685650,
  685650, 685680,
  685680, 685711,
  685711, 685741,
  685741, 685772,
  685772, 685803,
  685803, 685833,
  685833, 685864,
  685864, 685894,
  685894, 685925,
  685925, 685956,
  685956, 685984,
  685984, 686015,
  686015, 686045,
  686045, 686076,
  686076, 686106,
  686106, 686137,
  686137, 686168,
  686168, 686198,
  686198, 686229,
  686229, 686259,
  686259, 686290,
  686290, 686321,
  686321, 686350,
  686350, 686381,
  686381, 686411,
  686411, 686442,
  686442, 686472,
  686472, 686503,
  686503, 686534,
  686534, 686564,
  686564, 686595,
  686595, 686625,
  686625, 686656,
  686656, 686687,
  686687, 686715,
  686715, 686746,
  686746, 686776,
  686776, 686807,
  686807, 686837,
  686837, 686868,
  686868, 686899,
  686899, 686929,
  686929, 686960,
  686960, 686990,
  686990, 687021,
  687021, 687052,
  687052, 687080,
  687080, 687111,
  687111, 687141,
  687141, 687172,
  687172, 687202,
  687202, 687233,
  687233, 687264,
  687264, 687294,
  687294, 687325,
  687325, 687355,
  687355, 687386,
  687386, 687417,
  687417, 687445,
  687445, 687476,
  687476, 687506,
  687506, 687537,
  687537, 687567,
  687567, 687598,
  687598, 687629,
  687629, 687659,
  687659, 687690,
  687690, 687720,
  687720, 687751,
  687751, 687782,
  687782, 687811,
  687811, 687842,
  687842, 687872,
  687872, 687903,
  687903, 687933,
  687933, 687964,
  687964, 687995,
  687995, 688025,
  688025, 688056,
  688056, 688086,
  688086, 688117,
  688117, 688148,
  688148, 688176,
  688176, 688207,
  688207, 688237,
  688237, 688268,
  688268, 688298,
  688298, 688329,
  688329, 688360,
  688360, 688390,
  688390, 688421,
  688421, 688451,
  688451, 688482,
  688482, 688513,
  688513, 688541,
  688541, 688572,
  688572, 688602,
  688602, 688633,
  688633, 688663,
  688663, 688694,
  688694, 688725,
  688725, 688755,
  688755, 688786,
  688786, 688816,
  688816, 688847,
  688847, 688878,
  688878, 688906,
  688906, 688937,
  688937, 688967,
  688967, 688998,
  688998, 689028,
  689028, 689059,
  689059, 689090,
  689090, 689120,
  689120, 689151,
  689151, 689181,
  689181, 689212,
  689212, 689243,
  689243, 689272,
  689272, 689303,
  689303, 689333,
  689333, 689364,
  689364, 689394,
  689394, 689425,
  689425, 689456,
  689456, 689486,
  689486, 689517,
  689517, 689547,
  689547, 689578,
  689578, 689609,
  689609, 689637,
  689637, 689668,
  689668, 689698,
  689698, 689729,
  689729, 689759,
  689759, 689790,
  689790, 689821,
  689821, 689851,
  689851, 689882,
  689882, 689912,
  689912, 689943,
  689943, 689974,
  689974, 690002,
  690002, 690033,
  690033, 690063,
  690063, 690094,
  690094, 690124,
  690124, 690155,
  690155, 690186,
  690186, 690216,
  690216, 690247,
  690247, 690277,
  690277, 690308,
  690308, 690339,
  690339, 690367,
  690367, 690398,
  690398, 690428,
  690428, 690459,
  690459, 690489,
  690489, 690520,
  690520, 690551,
  690551, 690581,
  690581, 690612,
  690612, 690642,
  690642, 690673,
  690673, 690704,
  690704, 690733,
  690733, 690764,
  690764, 690794,
  690794, 690825,
  690825, 690855,
  690855, 690886,
  690886, 690917,
  690917, 690947,
  690947, 690978,
  690978, 691008,
  691008, 691039,
  691039, 691070,
  691070, 691098,
  691098, 691129,
  691129, 691159,
  691159, 691190,
  691190, 691220,
  691220, 691251,
  691251, 691282,
  691282, 691312,
  691312, 691343,
  691343, 691373,
  691373, 691404,
  691404, 691435,
  691435, 691463,
  691463, 691494,
  691494, 691524,
  691524, 691555,
  691555, 691585,
  691585, 691616,
  691616, 691647,
  691647, 691677,
  691677, 691708,
  691708, 691738,
  691738, 691769,
  691769, 691800,
  691800, 691828,
  691828, 691859,
  691859, 691889,
  691889, 691920,
  691920, 691950,
  691950, 691981,
  691981, 692012,
  692012, 692042,
  692042, 692073,
  692073, 692103,
  692103, 692134,
  692134, 692165,
  692165, 692194,
  692194, 692225,
  692225, 692255,
  692255, 692286,
  692286, 692316,
  692316, 692347,
  692347, 692378,
  692378, 692408,
  692408, 692439,
  692439, 692469,
  692469, 692500,
  692500, 692531,
  692531, 692559,
  692559, 692590,
  692590, 692620,
  692620, 692651,
  692651, 692681,
  692681, 692712,
  692712, 692743,
  692743, 692773,
  692773, 692804,
  692804, 692834,
  692834, 692865,
  692865, 692896,
  692896, 692924,
  692924, 692955,
  692955, 692985,
  692985, 693016,
  693016, 693046,
  693046, 693077,
  693077, 693108,
  693108, 693138,
  693138, 693169,
  693169, 693199,
  693199, 693230,
  693230, 693261,
  693261, 693289,
  693289, 693320,
  693320, 693350,
  693350, 693381,
  693381, 693411,
  693411, 693442,
  693442, 693473,
  693473, 693503,
  693503, 693534,
  693534, 693564,
  693564, 693595,
  693595, 693626,
  693626, 693654,
  693654, 693685,
  693685, 693715,
  693715, 693746,
  693746, 693776,
  693776, 693807,
  693807, 693838,
  693838, 693868,
  693868, 693899,
  693899, 693929,
  693929, 693960,
  693960, 693991,
  693991, 694019,
  694019, 694050,
  694050, 694080,
  694080, 694111,
  694111, 694141,
  694141, 694172,
  694172, 694203,
  694203, 694233,
  694233, 694264,
  694264, 694294,
  694294, 694325,
  694325, 694356,
  694356, 694384,
  694384, 694415,
  694415, 694445,
  694445, 694476,
  694476, 694506,
  694506, 694537,
  694537, 694568,
  694568, 694598,
  694598, 694629,
  694629, 694659,
  694659, 694690,
  694690, 694721,
  694721, 694749,
  694749, 694780,
  694780, 694810,
  694810, 694841,
  694841, 694871,
  694871, 694902,
  694902, 694933,
  694933, 694963,
  694963, 694994,
  694994, 695024,
  695024, 695055,
  695055, 695086,
  695086, 695115,
  695115, 695146,
  695146, 695176,
  695176, 695207,
  695207, 695237,
  695237, 695268,
  695268, 695299,
  695299, 695329,
  695329, 695360,
  695360, 695390,
  695390, 695421,
  695421, 695452,
  695452, 695480,
  695480, 695511,
  695511, 695541,
  695541, 695572,
  695572, 695602,
  695602, 695633,
  695633, 695664,
  695664, 695694,
  695694, 695725,
  695725, 695755,
  695755, 695786,
  695786, 695817,
  695817, 695845,
  695845, 695876,
  695876, 695906,
  695906, 695937,
  695937, 695967,
  695967, 695998,
  695998, 696029,
  696029, 696059,
  696059, 696090,
  696090, 696120,
  696120, 696151,
  696151, 696182,
  696182, 696210,
  696210, 696241,
  696241, 696271,
  696271, 696302,
  696302, 696332,
  696332, 696363,
  696363, 696394,
  696394, 696424,
  696424, 696455,
  696455, 696485,
  696485, 696516,
  696516, 696547,
  696547, 696576,
  696576, 696607,
  696607, 696637,
  696637, 696668,
  696668, 696698,
  696698, 696729,
  696729, 696760,
  696760, 696790,
  696790, 696821,
  696821, 696851,
  696851, 696882,
  696882, 696913,
  696913, 696941,
  696941, 696972,
  696972, 697002,
  697002, 697033,
  697033, 697063,
  697063, 697094,
  697094, 697125,
  697125, 697155,
  697155, 697186,
  697186, 697216,
  697216, 697247,
  697247, 697278,
  697278, 697306,
  697306, 697337,
  697337, 697367,
  697367, 697398,
  697398, 697428,
  697428, 697459,
  697459, 697490,
  697490, 697520,
  697520, 697551,
  697551, 697581,
  697581, 697612,
  697612, 697643,
  697643, 697671,
  697671, 697702,
  697702, 697732,
  697732, 697763,
  697763, 697793,
  697793, 697824,
  697824, 697855,
  697855, 697885,
  697885, 697916,
  697916, 697946,
  697946, 697977,
  697977, 698008,
  698008, 698037,
  698037, 698068,
  698068, 698098,
  698098, 698129,
  698129, 698159,
  698159, 698190,
  698190, 698221,
  698221, 698251,
  698251, 698282,
  698282, 698312,
  698312, 698343,
  698343, 698374,
  698374, 698402,
  698402, 698433,
  698433, 698463,
  698463, 698494,
  698494, 698524,
  698524, 698555,
  698555, 698586,
  698586, 698616,
  698616, 698647,
  698647, 698677,
  698677, 698708,
  698708, 698739,
  698739, 698767,
  698767, 698798,
  698798, 698828,
  698828, 698859,
  698859, 698889,
  698889, 698920,
  698920, 698951,
  698951, 698981,
  698981, 699012,
  699012, 699042,
  699042, 699073,
  699073, 699104,
  699104, 699132,
  699132, 699163,
  699163, 699193,
  699193, 699224,
  699224, 699254,
  699254, 699285,
  699285, 699316,
  699316, 699346,
  699346, 699377,
  699377, 699407,
  699407, 699438,
  699438, 699469,
  699469, 699498,
  699498, 699529,
  699529, 699559,
  699559, 699590,
  699590, 699620,
  699620, 699651,
  699651, 699682,
  699682, 699712,
  699712, 699743,
  699743, 699773,
  699773, 699804,
  699804, 699835,
  699835, 699863,
  699863, 699894,
  699894, 699924,
  699924, 699955,
  699955, 699985,
  699985, 700016,
  700016, 700047,
  700047, 700077,
  700077, 700108,
  700108, 700138,
  700138, 700169,
  700169, 700200,
  700200, 700228,
  700228, 700259,
  700259, 700289,
  700289, 700320,
  700320, 700350,
  700350, 700381,
  700381, 700412,
  700412, 700442,
  700442, 700473,
  700473, 700503,
  700503, 700534,
  700534, 700565,
  700565, 700593,
  700593, 700624,
  700624, 700654,
  700654, 700685,
  700685, 700715,
  700715, 700746,
  700746, 700777,
  700777, 700807,
  700807, 700838,
  700838, 700868,
  700868, 700899,
  700899, 700930,
  700930, 700959,
  700959, 700990,
  700990, 701020,
  701020, 701051,
  701051, 701081,
  701081, 701112,
  701112, 701143,
  701143, 701173,
  701173, 701204,
  701204, 701234,
  701234, 701265,
  701265, 701296,
  701296, 701324,
  701324, 701355,
  701355, 701385,
  701385, 701416,
  701416, 701446,
  701446, 701477,
  701477, 701508,
  701508, 701538,
  701538, 701569,
  701569, 701599,
  701599, 701630,
  701630, 701661,
  701661, 701689,
  701689, 701720,
  701720, 701750,
  701750, 701781,
  701781, 701811,
  701811, 701842,
  701842, 701873,
  701873, 701903,
  701903, 701934,
  701934, 701964,
  701964, 701995,
  701995, 702026,
  702026, 702054,
  702054, 702085,
  702085, 702115,
  702115, 702146,
  702146, 702176,
  702176, 702207,
  702207, 702238,
  702238, 702268,
  702268, 702299,
  702299, 702329,
  702329, 702360,
  702360, 702391,
  702391, 702420,
  702420, 702451,
  702451, 702481,
  702481, 702512,
  702512, 702542,
  702542, 702573,
  702573, 702604,
  702604, 702634,
  702634, 702665,
  702665, 702695,
  702695, 702726,
  702726, 702757,
  702757, 702785,
  702785, 702816,
  702816, 702846,
  702846, 702877,
  702877, 702907,
  702907, 702938,
  702938, 702969,
  702969, 702999,
  702999, 703030,
  703030, 703060,
  703060, 703091,
  703091, 703122,
  703122, 703150,
  703150, 703181,
  703181, 703211,
  703211, 703242,
  703242, 703272,
  703272, 703303,
  703303, 703334,
  703334, 703364,
  703364, 703395,
  703395, 703425,
  703425, 703456,
  703456, 703487,
  703487, 703515,
  703515, 703546,
  703546, 703576,
  703576, 703607,
  703607, 703637,
  703637, 703668,
  703668, 703699,
  703699, 703729,
  703729, 703760,
  703760, 703790,
  703790, 703821,
  703821, 703852,
  703852, 703881,
  703881, 703912,
  703912, 703942,
  703942, 703973,
  703973, 704003,
  704003, 704034,
  704034, 704065,
  704065, 704095,
  704095, 704126,
  704126, 704156,
  704156, 704187,
  704187, 704218,
  704218, 704246,
  704246, 704277,
  704277, 704307,
  704307, 704338,
  704338, 704368,
  704368, 704399,
  704399, 704430,
  704430, 704460,
  704460, 704491,
  704491, 704521,
  704521, 704552,
  704552, 704583,
  704583, 704611,
  704611, 704642,
  704642, 704672,
  704672, 704703,
  704703, 704733,
  704733, 704764,
  704764, 704795,
  704795, 704825,
  704825, 704856,
  704856, 704886,
  704886, 704917,
  704917, 704948,
  704948, 704976,
  704976, 705007,
  705007, 705037,
  705037, 705068,
  705068, 705098,
  705098, 705129,
  705129, 705160,
  705160, 705190,
  705190, 705221,
  705221, 705251,
  705251, 705282,
  705282, 705313,
  705313, 705342,
  705342, 705373,
  705373, 705403,
  705403, 705434,
  705434, 705464,
  705464, 705495,
  705495, 705526,
  705526, 705556,
  705556, 705587,
  705587, 705617,
  705617, 705648,
  705648, 705679,
  705679, 705707,
  705707, 705738,
  705738, 705768,
  705768, 705799,
  705799, 705829,
  705829, 705860,
  705860, 705891,
  705891, 705921,
  705921, 705952,
  705952, 705982,
  705982, 706013,
  706013, 706044,
  706044, 706072,
  706072, 706103,
  706103, 706133,
  706133, 706164,
  706164, 706194,
  706194, 706225,
  706225, 706256,
  706256, 706286,
  706286, 706317,
  706317, 706347,
  706347, 706378,
  706378, 706409,
  706409, 706437,
  706437, 706468,
  706468, 706498,
  706498, 706529,
  706529, 706559,
  706559, 706590,
  706590, 706621,
  706621, 706651,
  706651, 706682,
  706682, 706712,
  706712, 706743,
  706743, 706774,
  706774, 706803,
  706803, 706834,
  706834, 706864,
  706864, 706895,
  706895, 706925,
  706925, 706956,
  706956, 706987,
  706987, 707017,
  707017, 707048,
  707048, 707078,
  707078, 707109,
  707109, 707140,
  707140, 707168,
  707168, 707199,
  707199, 707229,
  707229, 707260,
  707260, 707290,
  707290, 707321,
  707321, 707352,
  707352, 707382,
  707382, 707413,
  707413, 707443,
  707443, 707474,
  707474, 707505,
  707505, 707533,
  707533, 707564,
  707564, 707594,
  707594, 707625,
  707625, 707655,
  707655, 707686,
  707686, 707717,
  707717, 707747,
  707747, 707778,
  707778, 707808,
  707808, 707839,
  707839, 707870,
  707870, 707898,
  707898, 707929,
  707929, 707959,
  707959, 707990,
  707990, 708020,
  708020, 708051,
  708051, 708082,
  708082, 708112,
  708112, 708143,
  708143, 708173,
  708173, 708204,
  708204, 708235,
  708235, 708264,
  708264, 708295,
  708295, 708325,
  708325, 708356,
  708356, 708386,
  708386, 708417,
  708417, 708448,
  708448, 708478,
  708478, 708509,
  708509, 708539,
  708539, 708570,
  708570, 708601,
  708601, 708629,
  708629, 708660,
  708660, 708690,
  708690, 708721,
  708721, 708751,
  708751, 708782,
  708782, 708813,
  708813, 708843,
  708843, 708874,
  708874, 708904,
  708904, 708935,
  708935, 708966,
  708966, 708994,
  708994, 709025,
  709025, 709055,
  709055, 709086,
  709086, 709116,
  709116, 709147,
  709147, 709178,
  709178, 709208,
  709208, 709239,
  709239, 709269,
  709269, 709300,
  709300, 709331,
  709331, 709359,
  709359, 709390,
  709390, 709420,
  709420, 709451,
  709451, 709481,
  709481, 709512,
  709512, 709543,
  709543, 709573,
  709573, 709604,
  709604, 709634,
  709634, 709665,
  709665, 709696,
  709696, 709725,
  709725, 709756,
  709756, 709786,
  709786, 709817,
  709817, 709847,
  709847, 709878,
  709878, 709909,
  709909, 709939,
  709939, 709970,
  709970, 710000,
  710000, 710031,
  710031, 710062,
  710062, 710090,
  710090, 710121,
  710121, 710151,
  710151, 710182,
  710182, 710212,
  710212, 710243,
  710243, 710274,
  710274, 710304,
  710304, 710335,
  710335, 710365,
  710365, 710396,
  710396, 710427,
  710427, 710455,
  710455, 710486,
  710486, 710516,
  710516, 710547,
  710547, 710577,
  710577, 710608,
  710608, 710639,
  710639, 710669,
  710669, 710700,
  710700, 710730,
  710730, 710761,
  710761, 710792,
  710792, 710820,
  710820, 710851,
  710851, 710881,
  710881, 710912,
  710912, 710942,
  710942, 710973,
  710973, 711004,
  711004, 711034,
  711034, 711065,
  711065, 711095,
  711095, 711126,
  711126, 711157,
  711157, 711186,
  711186, 711217,
  711217, 711247,
  711247, 711278,
  711278, 711308,
  711308, 711339,
  711339, 711370,
  711370, 711400,
  711400, 711431,
  711431, 711461,
  711461, 711492,
  711492, 711523,
  711523, 711551,
  711551, 711582,
  711582, 711612,
  711612, 711643,
  711643, 711673,
  711673, 711704,
  711704, 711735,
  711735, 711765,
  711765, 711796,
  711796, 711826,
  711826, 711857,
  711857, 711888,
  711888, 711916,
  711916, 711947,
  711947, 711977,
  711977, 712008,
  712008, 712038,
  712038, 712069,
  712069, 712100,
  712100, 712130,
  712130, 712161,
  712161, 712191,
  712191, 712222,
  712222, 712253,
  712253, 712281,
  712281, 712312,
  712312, 712342,
  712342, 712373,
  712373, 712403,
  712403, 712434,
  712434, 712465,
  712465, 712495,
  712495, 712526,
  712526, 712556,
  712556, 712587,
  712587, 712618,
  712618, 712647,
  712647, 712678,
  712678, 712708,
  712708, 712739,
  712739, 712769,
  712769, 712800,
  712800, 712831,
  712831, 712861,
  712861, 712892,
  712892, 712922,
  712922, 712953,
  712953, 712984,
  712984, 713012,
  713012, 713043,
  713043, 713073,
  713073, 713104,
  713104, 713134,
  713134, 713165,
  713165, 713196,
  713196, 713226,
  713226, 713257,
  713257, 713287,
  713287, 713318,
  713318, 713349,
  713349, 713377,
  713377, 713408,
  713408, 713438,
  713438, 713469,
  713469, 713499,
  713499, 713530,
  713530, 713561,
  713561, 713591,
  713591, 713622,
  713622, 713652,
  713652, 713683,
  713683, 713714,
  713714, 713742,
  713742, 713773,
  713773, 713803,
  713803, 713834,
  713834, 713864,
  713864, 713895,
  713895, 713926,
  713926, 713956,
  713956, 713987,
  713987, 714017,
  714017, 714048,
  714048, 714079,
  714079, 714108,
  714108, 714139,
  714139, 714169,
  714169, 714200,
  714200, 714230,
  714230, 714261,
  714261, 714292,
  714292, 714322,
  714322, 714353,
  714353, 714383,
  714383, 714414,
  714414, 714445,
  714445, 714473,
  714473, 714504,
  714504, 714534,
  714534, 714565,
  714565, 714595,
  714595, 714626,
  714626, 714657,
  714657, 714687,
  714687, 714718,
  714718, 714748,
  714748, 714779,
  714779, 714810,
  714810, 714838,
  714838, 714869,
  714869, 714899,
  714899, 714930,
  714930, 714960,
  714960, 714991,
  714991, 715022,
  715022, 715052,
  715052, 715083,
  715083, 715113,
  715113, 715144,
  715144, 715175,
  715175, 715203,
  715203, 715234,
  715234, 715264,
  715264, 715295,
  715295, 715325,
  715325, 715356,
  715356, 715387,
  715387, 715417,
  715417, 715448,
  715448, 715478,
  715478, 715509,
  715509, 715540,
  715540, 715569,
  715569, 715600,
  715600, 715630,
  715630, 715661,
  715661, 715691,
  715691, 715722,
  715722, 715753,
  715753, 715783,
  715783, 715814,
  715814, 715844,
  715844, 715875,
  715875, 715906,
  715906, 715934,
  715934, 715965,
  715965, 715995,
  715995, 716026,
  716026, 716056,
  716056, 716087,
  716087, 716118,
  716118, 716148,
  716148, 716179,
  716179, 716209,
  716209, 716240,
  716240, 716271,
  716271, 716299,
  716299, 716330,
  716330, 716360,
  716360, 716391,
  716391, 716421,
  716421, 716452,
  716452, 716483,
  716483, 716513,
  716513, 716544,
  716544, 716574,
  716574, 716605,
  716605, 716636,
  716636, 716664,
  716664, 716695,
  716695, 716725,
  716725, 716756,
  716756, 716786,
  716786, 716817,
  716817, 716848,
  716848, 716878,
  716878, 716909,
  716909, 716939,
  716939, 716970,
  716970, 717001,
  717001, 717030,
  717030, 717061,
  717061, 717091,
  717091, 717122,
  717122, 717152,
  717152, 717183,
  717183, 717214,
  717214, 717244,
  717244, 717275,
  717275, 717305,
  717305, 717336,
  717336, 717367,
  717367, 717395,
  717395, 717426,
  717426, 717456,
  717456, 717487,
  717487, 717517,
  717517, 717548,
  717548, 717579,
  717579, 717609,
  717609, 717640,
  717640, 717670,
  717670, 717701,
  717701, 717732,
  717732, 717760,
  717760, 717791,
  717791, 717821,
  717821, 717852,
  717852, 717882,
  717882, 717913,
  717913, 717944,
  717944, 717974,
  717974, 718005,
  718005, 718035,
  718035, 718066,
  718066, 718097,
  718097, 718125,
  718125, 718156,
  718156, 718186,
  718186, 718217,
  718217, 718247,
  718247, 718278,
  718278, 718309,
  718309, 718339,
  718339, 718370,
  718370, 718400,
  718400, 718431,
  718431, 718462,
  718462, 718491,
  718491, 718522,
  718522, 718552,
  718552, 718583,
  718583, 718613,
  718613, 718644,
  718644, 718675,
  718675, 718705,
  718705, 718736,
  718736, 718766,
  718766, 718797,
  718797, 718828,
  718828, 718856,
  718856, 718887,
  718887, 718917,
  718917, 718948,
  718948, 718978,
  718978, 719009,
  719009, 719040,
  719040, 719070,
  719070, 719101,
  719101, 719131,
  719131, 719162,
  719162, 719193,
  719193, 719221,
  719221, 719252,
  719252, 719282,
  719282, 719313,
  719313, 719343,
  719343, 719374,
  719374, 719405,
  719405, 719435,
  719435, 719466,
  719466, 719496,
  719496, 719527,
  719527, 719558,
  719558, 719586,
  719586, 719617,
  719617, 719647,
  719647, 719678,
  719678, 719708,
  719708, 719739,
  719739, 719770,
  719770, 719800,
  719800, 719831,
  719831, 719861,
  719861, 719892,
  719892, 719923,
  719923, 719952,
  719952, 719983,
  719983, 720013,
  720013, 720044,
  720044, 720074,
  720074, 720105,
  720105, 720136,
  720136, 720166,
  720166, 720197,
  720197, 720227,
  720227, 720258,
  720258, 720289,
  720289, 720317,
  720317, 720348,
  720348, 720378,
  720378, 720409,
  720409, 720439,
  720439, 720470,
  720470, 720501,
  720501, 720531,
  720531, 720562,
  720562, 720592,
  720592, 720623,
  720623, 720654,
  720654, 720682,
  720682, 720713,
  720713, 720743,
  720743, 720774,
  720774, 720804,
  720804, 720835,
  720835, 720866,
  720866, 720896,
  720896, 720927,
  720927, 720957,
  720957, 720988,
  720988, 721019,
  721019, 721047,
  721047, 721078,
  721078, 721108,
  721108, 721139,
  721139, 721169,
  721169, 721200,
  721200, 721231,
  721231, 721261,
  721261, 721292,
  721292, 721322,
  721322, 721353,
  721353, 721384,
  721384, 721413,
  721413, 721444,
  721444, 721474,
  721474, 721505,
  721505, 721535,
  721535, 721566,
  721566, 721597,
  721597, 721627,
  721627, 721658,
  721658, 721688,
  721688, 721719,
  721719, 721750,
  721750, 721778,
  721778, 721809,
  721809, 721839,
  721839, 721870,
  721870, 721900,
  721900, 721931,
  721931, 721962,
  721962, 721992,
  721992, 722023,
  722023, 722053,
  722053, 722084,
  722084, 722115,
  722115, 722143,
  722143, 722174,
  722174, 722204,
  722204, 722235,
  722235, 722265,
  722265, 722296,
  722296, 722327,
  722327, 722357,
  722357, 722388,
  722388, 722418,
  722418, 722449,
  722449, 722480,
  722480, 722508,
  722508, 722539,
  722539, 722569,
  722569, 722600,
  722600, 722630,
  722630, 722661,
  722661, 722692,
  722692, 722722,
  722722, 722753,
  722753, 722783,
  722783, 722814,
  722814, 722845,
  722845, 722874,
  722874, 722905,
  722905, 722935,
  722935, 722966,
  722966, 722996,
  722996, 723027,
  723027, 723058,
  723058, 723088,
  723088, 723119,
  723119, 723149,
  723149, 723180,
  723180, 723211,
  723211, 723239,
  723239, 723270,
  723270, 723300,
  723300, 723331,
  723331, 723361,
  723361, 723392,
  723392, 723423,
  723423, 723453,
  723453, 723484,
  723484, 723514,
  723514, 723545,
  723545, 723576,
  723576, 723604,
  723604, 723635,
  723635, 723665,
  723665, 723696,
  723696, 723726,
  723726, 723757,
  723757, 723788,
  723788, 723818,
  723818, 723849,
  723849, 723879,
  723879, 723910,
  723910, 723941,
  723941, 723969,
  723969, 724000,
  724000, 724030,
  724030, 724061,
  724061, 724091,
  724091, 724122,
  724122, 724153,
  724153, 724183,
  724183, 724214,
  724214, 724244,
  724244, 724275,
  724275, 724306,
  724306, 724335,
  724335, 724366,
  724366, 724396,
  724396, 724427,
  724427, 724457,
  724457, 724488,
  724488, 724519,
  724519, 724549,
  724549, 724580,
  724580, 724610,
  724610, 724641,
  724641, 724672,
  724672, 724700,
  724700, 724731,
  724731, 724761,
  724761, 724792,
  724792, 724822,
  724822, 724853,
  724853, 724884,
  724884, 724914,
  724914, 724945,
  724945, 724975,
  724975, 725006,
  725006, 725037,
  725037, 725065,
  725065, 725096,
  725096, 725126,
  725126, 725157,
  725157, 725187,
  725187, 725218,
  725218, 725249,
  725249, 725279,
  725279, 725310,
  725310, 725340,
  725340, 725371,
  725371, 725402,
  725402, 725430,
  725430, 725461,
  725461, 725491,
  725491, 725522,
  725522, 725552,
  725552, 725583,
  725583, 725614,
  725614, 725644,
  725644, 725675,
  725675, 725705,
  725705, 725736,
  725736, 725767,
  725767, 725796,
  725796, 725827,
  725827, 725857,
  725857, 725888,
  725888, 725918,
  725918, 725949,
  725949, 725980,
  725980, 726010,
  726010, 726041,
  726041, 726071,
  726071, 726102,
  726102, 726133,
  726133, 726161,
  726161, 726192,
  726192, 726222,
  726222, 726253,
  726253, 726283,
  726283, 726314,
  726314, 726345,
  726345, 726375,
  726375, 726406,
  726406, 726436,
  726436, 726467,
  726467, 726498,
  726498, 726526,
  726526, 726557,
  726557, 726587,
  726587, 726618,
  726618, 726648,
  726648, 726679,
  726679, 726710,
  726710, 726740,
  726740, 726771,
  726771, 726801,
  726801, 726832,
  726832, 726863,
  726863, 726891,
  726891, 726922,
  726922, 726952,
  726952, 726983,
  726983, 727013,
  727013, 727044,
  727044, 727075,
  727075, 727105,
  727105, 727136,
  727136, 727166,
  727166, 727197,
  727197, 727228,
  727228, 727257,
  727257, 727288,
  727288, 727318,
  727318, 727349,
  727349, 727379,
  727379, 727410,
  727410, 727441,
  727441, 727471,
  727471, 727502,
  727502, 727532,
  727532, 727563,
  727563, 727594,
  727594, 727622,
  727622, 727653,
  727653, 727683,
  727683, 727714,
  727714, 727744,
  727744, 727775,
  727775, 727806,
  727806, 727836,
  727836, 727867,
  727867, 727897,
  727897, 727928,
  727928, 727959,
  727959, 727987,
  727987, 728018,
  728018, 728048,
  728048, 728079,
  728079, 728109,
  728109, 728140,
  728140, 728171,
  728171, 728201,
  728201, 728232,
  728232, 728262,
  728262, 728293,
  728293, 728324,
  728324, 728352,
  728352, 728383,
  728383, 728413,
  728413, 728444,
  728444, 728474,
  728474, 728505,
  728505, 728536,
  728536, 728566,
  728566, 728597,
  728597, 728627,
  728627, 728658,
  728658, 728689,
  728689, 728718,
  728718, 728749,
  728749, 728779,
  728779, 728810,
  728810, 728840,
  728840, 728871,
  728871, 728902,
  728902, 728932,
  728932, 728963,
  728963, 728993,
  728993, 729024,
  729024, 729055,
  729055, 729083,
  729083, 729114,
  729114, 729144,
  729144, 729175,
  729175, 729205,
  729205, 729236,
  729236, 729267,
  729267, 729297,
  729297, 729328,
  729328, 729358,
  729358, 729389,
  729389, 729420,
  729420, 729448,
  729448, 729479,
  729479, 729509,
  729509, 729540,
  729540, 729570,
  729570, 729601,
  729601, 729632,
  729632, 729662,
  729662, 729693,
  729693, 729723,
  729723, 729754,
  729754, 729785,
  729785, 729813,
  729813, 729844,
  729844, 729874,
  729874, 729905,
  729905, 729935,
  729935, 729966,
  729966, 729997,
  729997, 730027,
  730027, 730058,
  730058, 730088,
  730088, 730119,
  730119, 730150,
  730150, 730179,
  730179, 730210,
  730210, 730240,
  730240, 730271,
  730271, 730301,
  730301, 730332,
  730332, 730363,
  730363, 730393,
  730393, 730424,
  730424, 730454,
  730454, 730485,
  730485, 730516,
  730516, 730544,
  730544, 730575,
  730575, 730605,
  730605, 730636,
  730636, 730666,
  730666, 730697,
  730697, 730728,
  730728, 730758,
  730758, 730789,
  730789, 730819,
  730819, 730850,
  730850, 730881,
  730881, 730909,
  730909, 730940,
  730940, 730970,
  730970, 731001,
  731001, 731031,
  731031, 731062,
  731062, 731093,
  731093, 731123,
  731123, 731154,
  731154, 731184,
  731184, 731215,
  731215, 731246,
  731246, 731274,
  731274, 731305,
  731305, 731335,
  731335, 731366,
  731366, 731396,
  731396, 731427,
  731427, 731458,
  731458, 731488,
  731488, 731519,
  731519, 731549,
  731549, 731580,
  731580, 731611,
  731611, 731640,
  731640, 731671,
  731671, 731701,
  731701, 731732,
  731732, 731762,
  731762, 731793,
  731793, 731824,
  731824, 731854,
  731854, 731885,
  731885, 731915,
  731915, 731946,
  731946, 731977,
  731977, 732005,
  732005, 732036,
  732036, 732066,
  732066, 732097,
  732097, 732127,
  732127, 732158,
  732158, 732189,
  732189, 732219,
  732219, 732250,
  732250, 732280,
  732280, 732311 ;

 lat = _ ;

 lon = _ ;

 z = _ ;

 temperature =
  _, _,
  _, _,
  _, _,
  _, _ ;
}
