netcdf test_mon_365_day {
dimensions:
	time = UNLIMITED ;
	lat = 2 ;
	lon = 2 ;
    bnds = 2 ;
variables:
	double time(time) ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1850-1-1" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
	double time_bnds(time, bnds) ;
	float lat ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "Latitude" ;
	float lon ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "Longitude" ;
	float z ;
		z:standard_name = "depth" ;
		z:positive = "down" ;
		z:units = "m" ;
		z:long_name = "Depth below surface" ;
	float temperature(time, lat, lon) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "deg_C" ;
		temperature:long_name = "Seawater Temperature" ;
		temperature:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:variable_id = "temp-max" ;
		:scenario = "sres-a1b" ;
		:dataset_id = "ukcp18-land-prob-25km" ;
		:prob_type = "sample" ;
		:frequency = "mon" ;
data:

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319,
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684,
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5,
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5,
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626,
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5, 1840.5, 1870, 1899.5, 1930,
    1960.5, 1991, 2021.5, 2052.5, 2083, 2113.5, 2144, 2174.5, 2205.5, 2235,
    2264.5, 2295, 2325.5, 2356, 2386.5, 2417.5, 2448, 2478.5, 2509, 2539.5,
    2570.5, 2600, 2629.5, 2660, 2690.5, 2721, 2751.5, 2782.5, 2813, 2843.5,
    2874, 2904.5, 2935.5, 2965, 2994.5, 3025, 3055.5, 3086, 3116.5, 3147.5,
    3178, 3208.5, 3239, 3269.5, 3300.5, 3330, 3359.5, 3390, 3420.5, 3451,
    3481.5, 3512.5, 3543, 3573.5, 3604, 3634.5, 3665.5, 3695, 3724.5, 3755,
    3785.5, 3816, 3846.5, 3877.5, 3908, 3938.5, 3969, 3999.5, 4030.5, 4060,
    4089.5, 4120, 4150.5, 4181, 4211.5, 4242.5, 4273, 4303.5, 4334, 4364.5,
    4395.5, 4425, 4454.5, 4485, 4515.5, 4546, 4576.5, 4607.5, 4638, 4668.5,
    4699, 4729.5, 4760.5, 4790, 4819.5, 4850, 4880.5, 4911, 4941.5, 4972.5,
    5003, 5033.5, 5064, 5094.5, 5125.5, 5155, 5184.5, 5215, 5245.5, 5276,
    5306.5, 5337.5, 5368, 5398.5, 5429, 5459.5, 5490.5, 5520, 5549.5, 5580,
    5610.5, 5641, 5671.5, 5702.5, 5733, 5763.5, 5794, 5824.5, 5855.5, 5885,
    5914.5, 5945, 5975.5, 6006, 6036.5, 6067.5, 6098, 6128.5, 6159, 6189.5,
    6220.5, 6250, 6279.5, 6310, 6340.5, 6371, 6401.5, 6432.5, 6463, 6493.5,
    6524, 6554.5, 6585.5, 6615, 6644.5, 6675, 6705.5, 6736, 6766.5, 6797.5,
    6828, 6858.5, 6889, 6919.5, 6950.5, 6980, 7009.5, 7040, 7070.5, 7101,
    7131.5, 7162.5, 7193, 7223.5, 7254, 7284.5, 7315.5, 7345, 7374.5, 7405,
    7435.5, 7466, 7496.5, 7527.5, 7558, 7588.5, 7619, 7649.5, 7680.5, 7710,
    7739.5, 7770, 7800.5, 7831, 7861.5, 7892.5, 7923, 7953.5, 7984, 8014.5,
    8045.5, 8075, 8104.5, 8135, 8165.5, 8196, 8226.5, 8257.5, 8288, 8318.5,
    8349, 8379.5, 8410.5, 8440, 8469.5, 8500, 8530.5, 8561, 8591.5, 8622.5,
    8653, 8683.5, 8714, 8744.5, 8775.5, 8805, 8834.5, 8865, 8895.5, 8926,
    8956.5, 8987.5, 9018, 9048.5, 9079, 9109.5, 9140.5, 9170, 9199.5, 9230,
    9260.5, 9291, 9321.5, 9352.5, 9383, 9413.5, 9444, 9474.5, 9505.5, 9535,
    9564.5, 9595, 9625.5, 9656, 9686.5, 9717.5, 9748, 9778.5, 9809, 9839.5,
    9870.5, 9900, 9929.5, 9960, 9990.5, 10021, 10051.5, 10082.5, 10113,
    10143.5, 10174, 10204.5, 10235.5, 10265, 10294.5, 10325, 10355.5, 10386,
    10416.5, 10447.5, 10478, 10508.5, 10539, 10569.5, 10600.5, 10630,
    10659.5, 10690, 10720.5, 10751, 10781.5, 10812.5, 10843, 10873.5, 10904,
    10934.5, 10965.5, 10995, 11024.5, 11055, 11085.5, 11116, 11146.5,
    11177.5, 11208, 11238.5, 11269, 11299.5, 11330.5, 11360, 11389.5, 11420,
    11450.5, 11481, 11511.5, 11542.5, 11573, 11603.5, 11634, 11664.5,
    11695.5, 11725, 11754.5, 11785, 11815.5, 11846, 11876.5, 11907.5, 11938,
    11968.5, 11999, 12029.5, 12060.5, 12090, 12119.5, 12150, 12180.5, 12211,
    12241.5, 12272.5, 12303, 12333.5, 12364, 12394.5, 12425.5, 12455,
    12484.5, 12515, 12545.5, 12576, 12606.5, 12637.5, 12668, 12698.5, 12729,
    12759.5, 12790.5, 12820, 12849.5, 12880, 12910.5, 12941, 12971.5,
    13002.5, 13033, 13063.5, 13094, 13124.5, 13155.5, 13185, 13214.5, 13245,
    13275.5, 13306, 13336.5, 13367.5, 13398, 13428.5, 13459, 13489.5,
    13520.5, 13550, 13579.5, 13610, 13640.5, 13671, 13701.5, 13732.5, 13763,
    13793.5, 13824, 13854.5, 13885.5, 13915, 13944.5, 13975, 14005.5, 14036,
    14066.5, 14097.5, 14128, 14158.5, 14189, 14219.5, 14250.5, 14280,
    14309.5, 14340, 14370.5, 14401, 14431.5, 14462.5, 14493, 14523.5, 14554,
    14584.5, 14615.5, 14645, 14674.5, 14705, 14735.5, 14766, 14796.5,
    14827.5, 14858, 14888.5, 14919, 14949.5, 14980.5, 15010, 15039.5, 15070,
    15100.5, 15131, 15161.5, 15192.5, 15223, 15253.5, 15284, 15314.5,
    15345.5, 15375, 15404.5, 15435, 15465.5, 15496, 15526.5, 15557.5, 15588,
    15618.5, 15649, 15679.5, 15710.5, 15740, 15769.5, 15800, 15830.5, 15861,
    15891.5, 15922.5, 15953, 15983.5, 16014, 16044.5, 16075.5, 16105,
    16134.5, 16165, 16195.5, 16226, 16256.5, 16287.5, 16318, 16348.5, 16379,
    16409.5, 16440.5, 16470, 16499.5, 16530, 16560.5, 16591, 16621.5,
    16652.5, 16683, 16713.5, 16744, 16774.5, 16805.5, 16835, 16864.5, 16895,
    16925.5, 16956, 16986.5, 17017.5, 17048, 17078.5, 17109, 17139.5,
    17170.5, 17200, 17229.5, 17260, 17290.5, 17321, 17351.5, 17382.5, 17413,
    17443.5, 17474, 17504.5, 17535.5, 17565, 17594.5, 17625, 17655.5, 17686,
    17716.5, 17747.5, 17778, 17808.5, 17839, 17869.5, 17900.5, 17930,
    17959.5, 17990, 18020.5, 18051, 18081.5, 18112.5, 18143, 18173.5, 18204,
    18234.5, 18265.5, 18295, 18324.5, 18355, 18385.5, 18416, 18446.5,
    18477.5, 18508, 18538.5, 18569, 18599.5, 18630.5, 18660, 18689.5, 18720,
    18750.5, 18781, 18811.5, 18842.5, 18873, 18903.5, 18934, 18964.5,
    18995.5, 19025, 19054.5, 19085, 19115.5, 19146, 19176.5, 19207.5, 19238,
    19268.5, 19299, 19329.5, 19360.5, 19390, 19419.5, 19450, 19480.5, 19511,
    19541.5, 19572.5, 19603, 19633.5, 19664, 19694.5, 19725.5, 19755,
    19784.5, 19815, 19845.5, 19876, 19906.5, 19937.5, 19968, 19998.5, 20029,
    20059.5, 20090.5, 20120, 20149.5, 20180, 20210.5, 20241, 20271.5,
    20302.5, 20333, 20363.5, 20394, 20424.5, 20455.5, 20485, 20514.5, 20545,
    20575.5, 20606, 20636.5, 20667.5, 20698, 20728.5, 20759, 20789.5,
    20820.5, 20850, 20879.5, 20910, 20940.5, 20971, 21001.5, 21032.5, 21063,
    21093.5, 21124, 21154.5, 21185.5, 21215, 21244.5, 21275, 21305.5, 21336,
    21366.5, 21397.5, 21428, 21458.5, 21489, 21519.5, 21550.5, 21580,
    21609.5, 21640, 21670.5, 21701, 21731.5, 21762.5, 21793, 21823.5, 21854,
    21884.5, 21915.5, 21945, 21974.5, 22005, 22035.5, 22066, 22096.5,
    22127.5, 22158, 22188.5, 22219, 22249.5, 22280.5, 22310, 22339.5, 22370,
    22400.5, 22431, 22461.5, 22492.5, 22523, 22553.5, 22584, 22614.5,
    22645.5, 22675, 22704.5, 22735, 22765.5, 22796, 22826.5, 22857.5, 22888,
    22918.5, 22949, 22979.5, 23010.5, 23040, 23069.5, 23100, 23130.5, 23161,
    23191.5, 23222.5, 23253, 23283.5, 23314, 23344.5, 23375.5, 23405,
    23434.5, 23465, 23495.5, 23526, 23556.5, 23587.5, 23618, 23648.5, 23679,
    23709.5, 23740.5, 23770, 23799.5, 23830, 23860.5, 23891, 23921.5,
    23952.5, 23983, 24013.5, 24044, 24074.5, 24105.5, 24135, 24164.5, 24195,
    24225.5, 24256, 24286.5, 24317.5, 24348, 24378.5, 24409, 24439.5,
    24470.5, 24500, 24529.5, 24560, 24590.5, 24621, 24651.5, 24682.5, 24713,
    24743.5, 24774, 24804.5, 24835.5, 24865, 24894.5, 24925, 24955.5, 24986,
    25016.5, 25047.5, 25078, 25108.5, 25139, 25169.5, 25200.5, 25230,
    25259.5, 25290, 25320.5, 25351, 25381.5, 25412.5, 25443, 25473.5, 25504,
    25534.5, 25565.5, 25595, 25624.5, 25655, 25685.5, 25716, 25746.5,
    25777.5, 25808, 25838.5, 25869, 25899.5, 25930.5, 25960, 25989.5, 26020,
    26050.5, 26081, 26111.5, 26142.5, 26173, 26203.5, 26234, 26264.5,
    26295.5, 26325, 26354.5, 26385, 26415.5, 26446, 26476.5, 26507.5, 26538,
    26568.5, 26599, 26629.5, 26660.5, 26690, 26719.5, 26750, 26780.5, 26811,
    26841.5, 26872.5, 26903, 26933.5, 26964, 26994.5, 27025.5, 27055,
    27084.5, 27115, 27145.5, 27176, 27206.5, 27237.5, 27268, 27298.5, 27329,
    27359.5, 27390.5, 27420, 27449.5, 27480, 27510.5, 27541, 27571.5,
    27602.5, 27633, 27663.5, 27694, 27724.5, 27755.5, 27785, 27814.5, 27845,
    27875.5, 27906, 27936.5, 27967.5, 27998, 28028.5, 28059, 28089.5,
    28120.5, 28150, 28179.5, 28210, 28240.5, 28271, 28301.5, 28332.5, 28363,
    28393.5, 28424, 28454.5, 28485.5, 28515, 28544.5, 28575, 28605.5, 28636,
    28666.5, 28697.5, 28728, 28758.5, 28789, 28819.5, 28850.5, 28880,
    28909.5, 28940, 28970.5, 29001, 29031.5, 29062.5, 29093, 29123.5, 29154,
    29184.5, 29215.5, 29245, 29274.5, 29305, 29335.5, 29366, 29396.5,
    29427.5, 29458, 29488.5, 29519, 29549.5, 29580.5, 29610, 29639.5, 29670,
    29700.5, 29731, 29761.5, 29792.5, 29823, 29853.5, 29884, 29914.5,
    29945.5, 29975, 30004.5, 30035, 30065.5, 30096, 30126.5, 30157.5, 30188,
    30218.5, 30249, 30279.5, 30310.5, 30340, 30369.5, 30400, 30430.5, 30461,
    30491.5, 30522.5, 30553, 30583.5, 30614, 30644.5, 30675.5, 30705,
    30734.5, 30765, 30795.5, 30826, 30856.5, 30887.5, 30918, 30948.5, 30979,
    31009.5, 31040.5, 31070, 31099.5, 31130, 31160.5, 31191, 31221.5,
    31252.5, 31283, 31313.5, 31344, 31374.5, 31405.5, 31435, 31464.5, 31495,
    31525.5, 31556, 31586.5, 31617.5, 31648, 31678.5, 31709, 31739.5,
    31770.5, 31800, 31829.5, 31860, 31890.5, 31921, 31951.5, 31982.5, 32013,
    32043.5, 32074, 32104.5, 32135.5, 32165, 32194.5, 32225, 32255.5, 32286,
    32316.5, 32347.5, 32378, 32408.5, 32439, 32469.5, 32500.5, 32530,
    32559.5, 32590, 32620.5, 32651, 32681.5, 32712.5, 32743, 32773.5, 32804,
    32834.5, 32865.5, 32895, 32924.5, 32955, 32985.5, 33016, 33046.5,
    33077.5, 33108, 33138.5, 33169, 33199.5, 33230.5, 33260, 33289.5, 33320,
    33350.5, 33381, 33411.5, 33442.5, 33473, 33503.5, 33534, 33564.5,
    33595.5, 33625, 33654.5, 33685, 33715.5, 33746, 33776.5, 33807.5, 33838,
    33868.5, 33899, 33929.5, 33960.5, 33990, 34019.5, 34050, 34080.5, 34111,
    34141.5, 34172.5, 34203, 34233.5, 34264, 34294.5, 34325.5, 34355,
    34384.5, 34415, 34445.5, 34476, 34506.5, 34537.5, 34568, 34598.5, 34629,
    34659.5, 34690.5, 34720, 34749.5, 34780, 34810.5, 34841, 34871.5,
    34902.5, 34933, 34963.5, 34994, 35024.5, 35055.5, 35085, 35114.5, 35145,
    35175.5, 35206, 35236.5, 35267.5, 35298, 35328.5, 35359, 35389.5,
    35420.5, 35450, 35479.5, 35510, 35540.5, 35571, 35601.5, 35632.5, 35663,
    35693.5, 35724, 35754.5, 35785.5, 35815, 35844.5, 35875, 35905.5, 35936,
    35966.5, 35997.5, 36028, 36058.5, 36089, 36119.5, 36150.5, 36180,
    36209.5, 36240, 36270.5, 36301, 36331.5, 36362.5, 36393, 36423.5, 36454,
    36484.5, 36515.5, 36545, 36574.5, 36605, 36635.5, 36666, 36696.5,
    36727.5, 36758, 36788.5, 36819, 36849.5, 36880.5, 36910, 36939.5, 36970,
    37000.5, 37031, 37061.5, 37092.5, 37123, 37153.5, 37184, 37214.5,
    37245.5, 37275, 37304.5, 37335, 37365.5, 37396, 37426.5, 37457.5, 37488,
    37518.5, 37549, 37579.5, 37610.5, 37640, 37669.5, 37700, 37730.5, 37761,
    37791.5, 37822.5, 37853, 37883.5, 37914, 37944.5, 37975.5, 38005,
    38034.5, 38065, 38095.5, 38126, 38156.5, 38187.5, 38218, 38248.5, 38279,
    38309.5, 38340.5, 38370, 38399.5, 38430, 38460.5, 38491, 38521.5,
    38552.5, 38583, 38613.5, 38644, 38674.5, 38705.5, 38735, 38764.5, 38795,
    38825.5, 38856, 38886.5, 38917.5, 38948, 38978.5, 39009, 39039.5,
    39070.5, 39100, 39129.5, 39160, 39190.5, 39221, 39251.5, 39282.5, 39313,
    39343.5, 39374, 39404.5, 39435.5, 39465, 39494.5, 39525, 39555.5, 39586,
    39616.5, 39647.5, 39678, 39708.5, 39739, 39769.5, 39800.5, 39830,
    39859.5, 39890, 39920.5, 39951, 39981.5, 40012.5, 40043, 40073.5, 40104,
    40134.5, 40165.5, 40195, 40224.5, 40255, 40285.5, 40316, 40346.5,
    40377.5, 40408, 40438.5, 40469, 40499.5, 40530.5, 40560, 40589.5, 40620,
    40650.5, 40681, 40711.5, 40742.5, 40773, 40803.5, 40834, 40864.5,
    40895.5, 40925, 40954.5, 40985, 41015.5, 41046, 41076.5, 41107.5, 41138,
    41168.5, 41199, 41229.5, 41260.5, 41290, 41319.5, 41350, 41380.5, 41411,
    41441.5, 41472.5, 41503, 41533.5, 41564, 41594.5, 41625.5, 41655,
    41684.5, 41715, 41745.5, 41776, 41806.5, 41837.5, 41868, 41898.5, 41929,
    41959.5, 41990.5, 42020, 42049.5, 42080, 42110.5, 42141, 42171.5,
    42202.5, 42233, 42263.5, 42294, 42324.5, 42355.5, 42385, 42414.5, 42445,
    42475.5, 42506, 42536.5, 42567.5, 42598, 42628.5, 42659, 42689.5,
    42720.5, 42750, 42779.5, 42810, 42840.5, 42871, 42901.5, 42932.5, 42963,
    42993.5, 43024, 43054.5, 43085.5, 43115, 43144.5, 43175, 43205.5, 43236,
    43266.5, 43297.5, 43328, 43358.5, 43389, 43419.5, 43450.5, 43480,
    43509.5, 43540, 43570.5, 43601, 43631.5, 43662.5, 43693, 43723.5, 43754,
    43784.5, 43815.5, 43845, 43874.5, 43905, 43935.5, 43966, 43996.5,
    44027.5, 44058, 44088.5, 44119, 44149.5, 44180.5, 44210, 44239.5, 44270,
    44300.5, 44331, 44361.5, 44392.5, 44423, 44453.5, 44484, 44514.5,
    44545.5, 44575, 44604.5, 44635, 44665.5, 44696, 44726.5, 44757.5, 44788,
    44818.5, 44849, 44879.5, 44910.5, 44940, 44969.5, 45000, 45030.5, 45061,
    45091.5, 45122.5, 45153, 45183.5, 45214, 45244.5, 45275.5, 45305,
    45334.5, 45365, 45395.5, 45426, 45456.5, 45487.5, 45518, 45548.5, 45579,
    45609.5, 45640.5, 45670, 45699.5, 45730, 45760.5, 45791, 45821.5,
    45852.5, 45883, 45913.5, 45944, 45974.5, 46005.5, 46035, 46064.5, 46095,
    46125.5, 46156, 46186.5, 46217.5, 46248, 46278.5, 46309, 46339.5,
    46370.5, 46400, 46429.5, 46460, 46490.5, 46521, 46551.5, 46582.5, 46613,
    46643.5, 46674, 46704.5, 46735.5, 46765, 46794.5, 46825, 46855.5, 46886,
    46916.5, 46947.5, 46978, 47008.5, 47039, 47069.5, 47100.5, 47130,
    47159.5, 47190, 47220.5, 47251, 47281.5, 47312.5, 47343, 47373.5, 47404,
    47434.5, 47465.5, 47495, 47524.5, 47555, 47585.5, 47616, 47646.5,
    47677.5, 47708, 47738.5, 47769, 47799.5, 47830.5, 47860, 47889.5, 47920,
    47950.5, 47981, 48011.5, 48042.5, 48073, 48103.5, 48134, 48164.5,
    48195.5, 48225, 48254.5, 48285, 48315.5, 48346, 48376.5, 48407.5, 48438,
    48468.5, 48499, 48529.5, 48560.5, 48590, 48619.5, 48650, 48680.5, 48711,
    48741.5, 48772.5, 48803, 48833.5, 48864, 48894.5, 48925.5, 48955,
    48984.5, 49015, 49045.5, 49076, 49106.5, 49137.5, 49168, 49198.5, 49229,
    49259.5, 49290.5, 49320, 49349.5, 49380, 49410.5, 49441, 49471.5,
    49502.5, 49533, 49563.5, 49594, 49624.5, 49655.5, 49685, 49714.5, 49745,
    49775.5, 49806, 49836.5, 49867.5, 49898, 49928.5, 49959, 49989.5,
    50020.5, 50050, 50079.5, 50110, 50140.5, 50171, 50201.5, 50232.5, 50263,
    50293.5, 50324, 50354.5, 50385.5, 50415, 50444.5, 50475, 50505.5, 50536,
    50566.5, 50597.5, 50628, 50658.5, 50689, 50719.5, 50750.5, 50780,
    50809.5, 50840, 50870.5, 50901, 50931.5, 50962.5, 50993, 51023.5, 51054,
    51084.5, 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5,
    51327.5, 51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570,
    51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5,
    51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 52088,
    52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 52330.5, 52361,
    52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 52575.5, 52605,
    52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 52818, 52848.5, 52879,
    52909.5, 52940.5, 52970, 52999.5, 53030, 53060.5, 53091, 53121.5,
    53152.5, 53183, 53213.5, 53244, 53274.5, 53305.5, 53335, 53364.5, 53395,
    53425.5, 53456, 53486.5, 53517.5, 53548, 53578.5, 53609, 53639.5,
    53670.5, 53700, 53729.5, 53760, 53790.5, 53821, 53851.5, 53882.5, 53913,
    53943.5, 53974, 54004.5, 54035.5, 54065, 54094.5, 54125, 54155.5, 54186,
    54216.5, 54247.5, 54278, 54308.5, 54339, 54369.5, 54400.5, 54430,
    54459.5, 54490, 54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704,
    54734.5, 54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5,
    54977.5, 55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220,
    55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5,
    55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 55738,
    55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 55980.5, 56011,
    56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 56225.5, 56255,
    56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 56468, 56498.5, 56529,
    56559.5, 56590.5, 56620, 56649.5, 56680, 56710.5, 56741, 56771.5,
    56802.5, 56833, 56863.5, 56894, 56924.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825,
  1825, 1856,
  1856, 1884,
  1884, 1915,
  1915, 1945,
  1945, 1976,
  1976, 2006,
  2006, 2037,
  2037, 2068,
  2068, 2098,
  2098, 2129,
  2129, 2159,
  2159, 2190,
  2190, 2221,
  2221, 2249,
  2249, 2280,
  2280, 2310,
  2310, 2341,
  2341, 2371,
  2371, 2402,
  2402, 2433,
  2433, 2463,
  2463, 2494,
  2494, 2524,
  2524, 2555,
  2555, 2586,
  2586, 2614,
  2614, 2645,
  2645, 2675,
  2675, 2706,
  2706, 2736,
  2736, 2767,
  2767, 2798,
  2798, 2828,
  2828, 2859,
  2859, 2889,
  2889, 2920,
  2920, 2951,
  2951, 2979,
  2979, 3010,
  3010, 3040,
  3040, 3071,
  3071, 3101,
  3101, 3132,
  3132, 3163,
  3163, 3193,
  3193, 3224,
  3224, 3254,
  3254, 3285,
  3285, 3316,
  3316, 3344,
  3344, 3375,
  3375, 3405,
  3405, 3436,
  3436, 3466,
  3466, 3497,
  3497, 3528,
  3528, 3558,
  3558, 3589,
  3589, 3619,
  3619, 3650,
  3650, 3681,
  3681, 3709,
  3709, 3740,
  3740, 3770,
  3770, 3801,
  3801, 3831,
  3831, 3862,
  3862, 3893,
  3893, 3923,
  3923, 3954,
  3954, 3984,
  3984, 4015,
  4015, 4046,
  4046, 4074,
  4074, 4105,
  4105, 4135,
  4135, 4166,
  4166, 4196,
  4196, 4227,
  4227, 4258,
  4258, 4288,
  4288, 4319,
  4319, 4349,
  4349, 4380,
  4380, 4411,
  4411, 4439,
  4439, 4470,
  4470, 4500,
  4500, 4531,
  4531, 4561,
  4561, 4592,
  4592, 4623,
  4623, 4653,
  4653, 4684,
  4684, 4714,
  4714, 4745,
  4745, 4776,
  4776, 4804,
  4804, 4835,
  4835, 4865,
  4865, 4896,
  4896, 4926,
  4926, 4957,
  4957, 4988,
  4988, 5018,
  5018, 5049,
  5049, 5079,
  5079, 5110,
  5110, 5141,
  5141, 5169,
  5169, 5200,
  5200, 5230,
  5230, 5261,
  5261, 5291,
  5291, 5322,
  5322, 5353,
  5353, 5383,
  5383, 5414,
  5414, 5444,
  5444, 5475,
  5475, 5506,
  5506, 5534,
  5534, 5565,
  5565, 5595,
  5595, 5626,
  5626, 5656,
  5656, 5687,
  5687, 5718,
  5718, 5748,
  5748, 5779,
  5779, 5809,
  5809, 5840,
  5840, 5871,
  5871, 5899,
  5899, 5930,
  5930, 5960,
  5960, 5991,
  5991, 6021,
  6021, 6052,
  6052, 6083,
  6083, 6113,
  6113, 6144,
  6144, 6174,
  6174, 6205,
  6205, 6236,
  6236, 6264,
  6264, 6295,
  6295, 6325,
  6325, 6356,
  6356, 6386,
  6386, 6417,
  6417, 6448,
  6448, 6478,
  6478, 6509,
  6509, 6539,
  6539, 6570,
  6570, 6601,
  6601, 6629,
  6629, 6660,
  6660, 6690,
  6690, 6721,
  6721, 6751,
  6751, 6782,
  6782, 6813,
  6813, 6843,
  6843, 6874,
  6874, 6904,
  6904, 6935,
  6935, 6966,
  6966, 6994,
  6994, 7025,
  7025, 7055,
  7055, 7086,
  7086, 7116,
  7116, 7147,
  7147, 7178,
  7178, 7208,
  7208, 7239,
  7239, 7269,
  7269, 7300,
  7300, 7331,
  7331, 7359,
  7359, 7390,
  7390, 7420,
  7420, 7451,
  7451, 7481,
  7481, 7512,
  7512, 7543,
  7543, 7573,
  7573, 7604,
  7604, 7634,
  7634, 7665,
  7665, 7696,
  7696, 7724,
  7724, 7755,
  7755, 7785,
  7785, 7816,
  7816, 7846,
  7846, 7877,
  7877, 7908,
  7908, 7938,
  7938, 7969,
  7969, 7999,
  7999, 8030,
  8030, 8061,
  8061, 8089,
  8089, 8120,
  8120, 8150,
  8150, 8181,
  8181, 8211,
  8211, 8242,
  8242, 8273,
  8273, 8303,
  8303, 8334,
  8334, 8364,
  8364, 8395,
  8395, 8426,
  8426, 8454,
  8454, 8485,
  8485, 8515,
  8515, 8546,
  8546, 8576,
  8576, 8607,
  8607, 8638,
  8638, 8668,
  8668, 8699,
  8699, 8729,
  8729, 8760,
  8760, 8791,
  8791, 8819,
  8819, 8850,
  8850, 8880,
  8880, 8911,
  8911, 8941,
  8941, 8972,
  8972, 9003,
  9003, 9033,
  9033, 9064,
  9064, 9094,
  9094, 9125,
  9125, 9156,
  9156, 9184,
  9184, 9215,
  9215, 9245,
  9245, 9276,
  9276, 9306,
  9306, 9337,
  9337, 9368,
  9368, 9398,
  9398, 9429,
  9429, 9459,
  9459, 9490,
  9490, 9521,
  9521, 9549,
  9549, 9580,
  9580, 9610,
  9610, 9641,
  9641, 9671,
  9671, 9702,
  9702, 9733,
  9733, 9763,
  9763, 9794,
  9794, 9824,
  9824, 9855,
  9855, 9886,
  9886, 9914,
  9914, 9945,
  9945, 9975,
  9975, 10006,
  10006, 10036,
  10036, 10067,
  10067, 10098,
  10098, 10128,
  10128, 10159,
  10159, 10189,
  10189, 10220,
  10220, 10251,
  10251, 10279,
  10279, 10310,
  10310, 10340,
  10340, 10371,
  10371, 10401,
  10401, 10432,
  10432, 10463,
  10463, 10493,
  10493, 10524,
  10524, 10554,
  10554, 10585,
  10585, 10616,
  10616, 10644,
  10644, 10675,
  10675, 10705,
  10705, 10736,
  10736, 10766,
  10766, 10797,
  10797, 10828,
  10828, 10858,
  10858, 10889,
  10889, 10919,
  10919, 10950,
  10950, 10981,
  10981, 11009,
  11009, 11040,
  11040, 11070,
  11070, 11101,
  11101, 11131,
  11131, 11162,
  11162, 11193,
  11193, 11223,
  11223, 11254,
  11254, 11284,
  11284, 11315,
  11315, 11346,
  11346, 11374,
  11374, 11405,
  11405, 11435,
  11435, 11466,
  11466, 11496,
  11496, 11527,
  11527, 11558,
  11558, 11588,
  11588, 11619,
  11619, 11649,
  11649, 11680,
  11680, 11711,
  11711, 11739,
  11739, 11770,
  11770, 11800,
  11800, 11831,
  11831, 11861,
  11861, 11892,
  11892, 11923,
  11923, 11953,
  11953, 11984,
  11984, 12014,
  12014, 12045,
  12045, 12076,
  12076, 12104,
  12104, 12135,
  12135, 12165,
  12165, 12196,
  12196, 12226,
  12226, 12257,
  12257, 12288,
  12288, 12318,
  12318, 12349,
  12349, 12379,
  12379, 12410,
  12410, 12441,
  12441, 12469,
  12469, 12500,
  12500, 12530,
  12530, 12561,
  12561, 12591,
  12591, 12622,
  12622, 12653,
  12653, 12683,
  12683, 12714,
  12714, 12744,
  12744, 12775,
  12775, 12806,
  12806, 12834,
  12834, 12865,
  12865, 12895,
  12895, 12926,
  12926, 12956,
  12956, 12987,
  12987, 13018,
  13018, 13048,
  13048, 13079,
  13079, 13109,
  13109, 13140,
  13140, 13171,
  13171, 13199,
  13199, 13230,
  13230, 13260,
  13260, 13291,
  13291, 13321,
  13321, 13352,
  13352, 13383,
  13383, 13413,
  13413, 13444,
  13444, 13474,
  13474, 13505,
  13505, 13536,
  13536, 13564,
  13564, 13595,
  13595, 13625,
  13625, 13656,
  13656, 13686,
  13686, 13717,
  13717, 13748,
  13748, 13778,
  13778, 13809,
  13809, 13839,
  13839, 13870,
  13870, 13901,
  13901, 13929,
  13929, 13960,
  13960, 13990,
  13990, 14021,
  14021, 14051,
  14051, 14082,
  14082, 14113,
  14113, 14143,
  14143, 14174,
  14174, 14204,
  14204, 14235,
  14235, 14266,
  14266, 14294,
  14294, 14325,
  14325, 14355,
  14355, 14386,
  14386, 14416,
  14416, 14447,
  14447, 14478,
  14478, 14508,
  14508, 14539,
  14539, 14569,
  14569, 14600,
  14600, 14631,
  14631, 14659,
  14659, 14690,
  14690, 14720,
  14720, 14751,
  14751, 14781,
  14781, 14812,
  14812, 14843,
  14843, 14873,
  14873, 14904,
  14904, 14934,
  14934, 14965,
  14965, 14996,
  14996, 15024,
  15024, 15055,
  15055, 15085,
  15085, 15116,
  15116, 15146,
  15146, 15177,
  15177, 15208,
  15208, 15238,
  15238, 15269,
  15269, 15299,
  15299, 15330,
  15330, 15361,
  15361, 15389,
  15389, 15420,
  15420, 15450,
  15450, 15481,
  15481, 15511,
  15511, 15542,
  15542, 15573,
  15573, 15603,
  15603, 15634,
  15634, 15664,
  15664, 15695,
  15695, 15726,
  15726, 15754,
  15754, 15785,
  15785, 15815,
  15815, 15846,
  15846, 15876,
  15876, 15907,
  15907, 15938,
  15938, 15968,
  15968, 15999,
  15999, 16029,
  16029, 16060,
  16060, 16091,
  16091, 16119,
  16119, 16150,
  16150, 16180,
  16180, 16211,
  16211, 16241,
  16241, 16272,
  16272, 16303,
  16303, 16333,
  16333, 16364,
  16364, 16394,
  16394, 16425,
  16425, 16456,
  16456, 16484,
  16484, 16515,
  16515, 16545,
  16545, 16576,
  16576, 16606,
  16606, 16637,
  16637, 16668,
  16668, 16698,
  16698, 16729,
  16729, 16759,
  16759, 16790,
  16790, 16821,
  16821, 16849,
  16849, 16880,
  16880, 16910,
  16910, 16941,
  16941, 16971,
  16971, 17002,
  17002, 17033,
  17033, 17063,
  17063, 17094,
  17094, 17124,
  17124, 17155,
  17155, 17186,
  17186, 17214,
  17214, 17245,
  17245, 17275,
  17275, 17306,
  17306, 17336,
  17336, 17367,
  17367, 17398,
  17398, 17428,
  17428, 17459,
  17459, 17489,
  17489, 17520,
  17520, 17551,
  17551, 17579,
  17579, 17610,
  17610, 17640,
  17640, 17671,
  17671, 17701,
  17701, 17732,
  17732, 17763,
  17763, 17793,
  17793, 17824,
  17824, 17854,
  17854, 17885,
  17885, 17916,
  17916, 17944,
  17944, 17975,
  17975, 18005,
  18005, 18036,
  18036, 18066,
  18066, 18097,
  18097, 18128,
  18128, 18158,
  18158, 18189,
  18189, 18219,
  18219, 18250,
  18250, 18281,
  18281, 18309,
  18309, 18340,
  18340, 18370,
  18370, 18401,
  18401, 18431,
  18431, 18462,
  18462, 18493,
  18493, 18523,
  18523, 18554,
  18554, 18584,
  18584, 18615,
  18615, 18646,
  18646, 18674,
  18674, 18705,
  18705, 18735,
  18735, 18766,
  18766, 18796,
  18796, 18827,
  18827, 18858,
  18858, 18888,
  18888, 18919,
  18919, 18949,
  18949, 18980,
  18980, 19011,
  19011, 19039,
  19039, 19070,
  19070, 19100,
  19100, 19131,
  19131, 19161,
  19161, 19192,
  19192, 19223,
  19223, 19253,
  19253, 19284,
  19284, 19314,
  19314, 19345,
  19345, 19376,
  19376, 19404,
  19404, 19435,
  19435, 19465,
  19465, 19496,
  19496, 19526,
  19526, 19557,
  19557, 19588,
  19588, 19618,
  19618, 19649,
  19649, 19679,
  19679, 19710,
  19710, 19741,
  19741, 19769,
  19769, 19800,
  19800, 19830,
  19830, 19861,
  19861, 19891,
  19891, 19922,
  19922, 19953,
  19953, 19983,
  19983, 20014,
  20014, 20044,
  20044, 20075,
  20075, 20106,
  20106, 20134,
  20134, 20165,
  20165, 20195,
  20195, 20226,
  20226, 20256,
  20256, 20287,
  20287, 20318,
  20318, 20348,
  20348, 20379,
  20379, 20409,
  20409, 20440,
  20440, 20471,
  20471, 20499,
  20499, 20530,
  20530, 20560,
  20560, 20591,
  20591, 20621,
  20621, 20652,
  20652, 20683,
  20683, 20713,
  20713, 20744,
  20744, 20774,
  20774, 20805,
  20805, 20836,
  20836, 20864,
  20864, 20895,
  20895, 20925,
  20925, 20956,
  20956, 20986,
  20986, 21017,
  21017, 21048,
  21048, 21078,
  21078, 21109,
  21109, 21139,
  21139, 21170,
  21170, 21201,
  21201, 21229,
  21229, 21260,
  21260, 21290,
  21290, 21321,
  21321, 21351,
  21351, 21382,
  21382, 21413,
  21413, 21443,
  21443, 21474,
  21474, 21504,
  21504, 21535,
  21535, 21566,
  21566, 21594,
  21594, 21625,
  21625, 21655,
  21655, 21686,
  21686, 21716,
  21716, 21747,
  21747, 21778,
  21778, 21808,
  21808, 21839,
  21839, 21869,
  21869, 21900,
  21900, 21931,
  21931, 21959,
  21959, 21990,
  21990, 22020,
  22020, 22051,
  22051, 22081,
  22081, 22112,
  22112, 22143,
  22143, 22173,
  22173, 22204,
  22204, 22234,
  22234, 22265,
  22265, 22296,
  22296, 22324,
  22324, 22355,
  22355, 22385,
  22385, 22416,
  22416, 22446,
  22446, 22477,
  22477, 22508,
  22508, 22538,
  22538, 22569,
  22569, 22599,
  22599, 22630,
  22630, 22661,
  22661, 22689,
  22689, 22720,
  22720, 22750,
  22750, 22781,
  22781, 22811,
  22811, 22842,
  22842, 22873,
  22873, 22903,
  22903, 22934,
  22934, 22964,
  22964, 22995,
  22995, 23026,
  23026, 23054,
  23054, 23085,
  23085, 23115,
  23115, 23146,
  23146, 23176,
  23176, 23207,
  23207, 23238,
  23238, 23268,
  23268, 23299,
  23299, 23329,
  23329, 23360,
  23360, 23391,
  23391, 23419,
  23419, 23450,
  23450, 23480,
  23480, 23511,
  23511, 23541,
  23541, 23572,
  23572, 23603,
  23603, 23633,
  23633, 23664,
  23664, 23694,
  23694, 23725,
  23725, 23756,
  23756, 23784,
  23784, 23815,
  23815, 23845,
  23845, 23876,
  23876, 23906,
  23906, 23937,
  23937, 23968,
  23968, 23998,
  23998, 24029,
  24029, 24059,
  24059, 24090,
  24090, 24121,
  24121, 24149,
  24149, 24180,
  24180, 24210,
  24210, 24241,
  24241, 24271,
  24271, 24302,
  24302, 24333,
  24333, 24363,
  24363, 24394,
  24394, 24424,
  24424, 24455,
  24455, 24486,
  24486, 24514,
  24514, 24545,
  24545, 24575,
  24575, 24606,
  24606, 24636,
  24636, 24667,
  24667, 24698,
  24698, 24728,
  24728, 24759,
  24759, 24789,
  24789, 24820,
  24820, 24851,
  24851, 24879,
  24879, 24910,
  24910, 24940,
  24940, 24971,
  24971, 25001,
  25001, 25032,
  25032, 25063,
  25063, 25093,
  25093, 25124,
  25124, 25154,
  25154, 25185,
  25185, 25216,
  25216, 25244,
  25244, 25275,
  25275, 25305,
  25305, 25336,
  25336, 25366,
  25366, 25397,
  25397, 25428,
  25428, 25458,
  25458, 25489,
  25489, 25519,
  25519, 25550,
  25550, 25581,
  25581, 25609,
  25609, 25640,
  25640, 25670,
  25670, 25701,
  25701, 25731,
  25731, 25762,
  25762, 25793,
  25793, 25823,
  25823, 25854,
  25854, 25884,
  25884, 25915,
  25915, 25946,
  25946, 25974,
  25974, 26005,
  26005, 26035,
  26035, 26066,
  26066, 26096,
  26096, 26127,
  26127, 26158,
  26158, 26188,
  26188, 26219,
  26219, 26249,
  26249, 26280,
  26280, 26311,
  26311, 26339,
  26339, 26370,
  26370, 26400,
  26400, 26431,
  26431, 26461,
  26461, 26492,
  26492, 26523,
  26523, 26553,
  26553, 26584,
  26584, 26614,
  26614, 26645,
  26645, 26676,
  26676, 26704,
  26704, 26735,
  26735, 26765,
  26765, 26796,
  26796, 26826,
  26826, 26857,
  26857, 26888,
  26888, 26918,
  26918, 26949,
  26949, 26979,
  26979, 27010,
  27010, 27041,
  27041, 27069,
  27069, 27100,
  27100, 27130,
  27130, 27161,
  27161, 27191,
  27191, 27222,
  27222, 27253,
  27253, 27283,
  27283, 27314,
  27314, 27344,
  27344, 27375,
  27375, 27406,
  27406, 27434,
  27434, 27465,
  27465, 27495,
  27495, 27526,
  27526, 27556,
  27556, 27587,
  27587, 27618,
  27618, 27648,
  27648, 27679,
  27679, 27709,
  27709, 27740,
  27740, 27771,
  27771, 27799,
  27799, 27830,
  27830, 27860,
  27860, 27891,
  27891, 27921,
  27921, 27952,
  27952, 27983,
  27983, 28013,
  28013, 28044,
  28044, 28074,
  28074, 28105,
  28105, 28136,
  28136, 28164,
  28164, 28195,
  28195, 28225,
  28225, 28256,
  28256, 28286,
  28286, 28317,
  28317, 28348,
  28348, 28378,
  28378, 28409,
  28409, 28439,
  28439, 28470,
  28470, 28501,
  28501, 28529,
  28529, 28560,
  28560, 28590,
  28590, 28621,
  28621, 28651,
  28651, 28682,
  28682, 28713,
  28713, 28743,
  28743, 28774,
  28774, 28804,
  28804, 28835,
  28835, 28866,
  28866, 28894,
  28894, 28925,
  28925, 28955,
  28955, 28986,
  28986, 29016,
  29016, 29047,
  29047, 29078,
  29078, 29108,
  29108, 29139,
  29139, 29169,
  29169, 29200,
  29200, 29231,
  29231, 29259,
  29259, 29290,
  29290, 29320,
  29320, 29351,
  29351, 29381,
  29381, 29412,
  29412, 29443,
  29443, 29473,
  29473, 29504,
  29504, 29534,
  29534, 29565,
  29565, 29596,
  29596, 29624,
  29624, 29655,
  29655, 29685,
  29685, 29716,
  29716, 29746,
  29746, 29777,
  29777, 29808,
  29808, 29838,
  29838, 29869,
  29869, 29899,
  29899, 29930,
  29930, 29961,
  29961, 29989,
  29989, 30020,
  30020, 30050,
  30050, 30081,
  30081, 30111,
  30111, 30142,
  30142, 30173,
  30173, 30203,
  30203, 30234,
  30234, 30264,
  30264, 30295,
  30295, 30326,
  30326, 30354,
  30354, 30385,
  30385, 30415,
  30415, 30446,
  30446, 30476,
  30476, 30507,
  30507, 30538,
  30538, 30568,
  30568, 30599,
  30599, 30629,
  30629, 30660,
  30660, 30691,
  30691, 30719,
  30719, 30750,
  30750, 30780,
  30780, 30811,
  30811, 30841,
  30841, 30872,
  30872, 30903,
  30903, 30933,
  30933, 30964,
  30964, 30994,
  30994, 31025,
  31025, 31056,
  31056, 31084,
  31084, 31115,
  31115, 31145,
  31145, 31176,
  31176, 31206,
  31206, 31237,
  31237, 31268,
  31268, 31298,
  31298, 31329,
  31329, 31359,
  31359, 31390,
  31390, 31421,
  31421, 31449,
  31449, 31480,
  31480, 31510,
  31510, 31541,
  31541, 31571,
  31571, 31602,
  31602, 31633,
  31633, 31663,
  31663, 31694,
  31694, 31724,
  31724, 31755,
  31755, 31786,
  31786, 31814,
  31814, 31845,
  31845, 31875,
  31875, 31906,
  31906, 31936,
  31936, 31967,
  31967, 31998,
  31998, 32028,
  32028, 32059,
  32059, 32089,
  32089, 32120,
  32120, 32151,
  32151, 32179,
  32179, 32210,
  32210, 32240,
  32240, 32271,
  32271, 32301,
  32301, 32332,
  32332, 32363,
  32363, 32393,
  32393, 32424,
  32424, 32454,
  32454, 32485,
  32485, 32516,
  32516, 32544,
  32544, 32575,
  32575, 32605,
  32605, 32636,
  32636, 32666,
  32666, 32697,
  32697, 32728,
  32728, 32758,
  32758, 32789,
  32789, 32819,
  32819, 32850,
  32850, 32881,
  32881, 32909,
  32909, 32940,
  32940, 32970,
  32970, 33001,
  33001, 33031,
  33031, 33062,
  33062, 33093,
  33093, 33123,
  33123, 33154,
  33154, 33184,
  33184, 33215,
  33215, 33246,
  33246, 33274,
  33274, 33305,
  33305, 33335,
  33335, 33366,
  33366, 33396,
  33396, 33427,
  33427, 33458,
  33458, 33488,
  33488, 33519,
  33519, 33549,
  33549, 33580,
  33580, 33611,
  33611, 33639,
  33639, 33670,
  33670, 33700,
  33700, 33731,
  33731, 33761,
  33761, 33792,
  33792, 33823,
  33823, 33853,
  33853, 33884,
  33884, 33914,
  33914, 33945,
  33945, 33976,
  33976, 34004,
  34004, 34035,
  34035, 34065,
  34065, 34096,
  34096, 34126,
  34126, 34157,
  34157, 34188,
  34188, 34218,
  34218, 34249,
  34249, 34279,
  34279, 34310,
  34310, 34341,
  34341, 34369,
  34369, 34400,
  34400, 34430,
  34430, 34461,
  34461, 34491,
  34491, 34522,
  34522, 34553,
  34553, 34583,
  34583, 34614,
  34614, 34644,
  34644, 34675,
  34675, 34706,
  34706, 34734,
  34734, 34765,
  34765, 34795,
  34795, 34826,
  34826, 34856,
  34856, 34887,
  34887, 34918,
  34918, 34948,
  34948, 34979,
  34979, 35009,
  35009, 35040,
  35040, 35071,
  35071, 35099,
  35099, 35130,
  35130, 35160,
  35160, 35191,
  35191, 35221,
  35221, 35252,
  35252, 35283,
  35283, 35313,
  35313, 35344,
  35344, 35374,
  35374, 35405,
  35405, 35436,
  35436, 35464,
  35464, 35495,
  35495, 35525,
  35525, 35556,
  35556, 35586,
  35586, 35617,
  35617, 35648,
  35648, 35678,
  35678, 35709,
  35709, 35739,
  35739, 35770,
  35770, 35801,
  35801, 35829,
  35829, 35860,
  35860, 35890,
  35890, 35921,
  35921, 35951,
  35951, 35982,
  35982, 36013,
  36013, 36043,
  36043, 36074,
  36074, 36104,
  36104, 36135,
  36135, 36166,
  36166, 36194,
  36194, 36225,
  36225, 36255,
  36255, 36286,
  36286, 36316,
  36316, 36347,
  36347, 36378,
  36378, 36408,
  36408, 36439,
  36439, 36469,
  36469, 36500,
  36500, 36531,
  36531, 36559,
  36559, 36590,
  36590, 36620,
  36620, 36651,
  36651, 36681,
  36681, 36712,
  36712, 36743,
  36743, 36773,
  36773, 36804,
  36804, 36834,
  36834, 36865,
  36865, 36896,
  36896, 36924,
  36924, 36955,
  36955, 36985,
  36985, 37016,
  37016, 37046,
  37046, 37077,
  37077, 37108,
  37108, 37138,
  37138, 37169,
  37169, 37199,
  37199, 37230,
  37230, 37261,
  37261, 37289,
  37289, 37320,
  37320, 37350,
  37350, 37381,
  37381, 37411,
  37411, 37442,
  37442, 37473,
  37473, 37503,
  37503, 37534,
  37534, 37564,
  37564, 37595,
  37595, 37626,
  37626, 37654,
  37654, 37685,
  37685, 37715,
  37715, 37746,
  37746, 37776,
  37776, 37807,
  37807, 37838,
  37838, 37868,
  37868, 37899,
  37899, 37929,
  37929, 37960,
  37960, 37991,
  37991, 38019,
  38019, 38050,
  38050, 38080,
  38080, 38111,
  38111, 38141,
  38141, 38172,
  38172, 38203,
  38203, 38233,
  38233, 38264,
  38264, 38294,
  38294, 38325,
  38325, 38356,
  38356, 38384,
  38384, 38415,
  38415, 38445,
  38445, 38476,
  38476, 38506,
  38506, 38537,
  38537, 38568,
  38568, 38598,
  38598, 38629,
  38629, 38659,
  38659, 38690,
  38690, 38721,
  38721, 38749,
  38749, 38780,
  38780, 38810,
  38810, 38841,
  38841, 38871,
  38871, 38902,
  38902, 38933,
  38933, 38963,
  38963, 38994,
  38994, 39024,
  39024, 39055,
  39055, 39086,
  39086, 39114,
  39114, 39145,
  39145, 39175,
  39175, 39206,
  39206, 39236,
  39236, 39267,
  39267, 39298,
  39298, 39328,
  39328, 39359,
  39359, 39389,
  39389, 39420,
  39420, 39451,
  39451, 39479,
  39479, 39510,
  39510, 39540,
  39540, 39571,
  39571, 39601,
  39601, 39632,
  39632, 39663,
  39663, 39693,
  39693, 39724,
  39724, 39754,
  39754, 39785,
  39785, 39816,
  39816, 39844,
  39844, 39875,
  39875, 39905,
  39905, 39936,
  39936, 39966,
  39966, 39997,
  39997, 40028,
  40028, 40058,
  40058, 40089,
  40089, 40119,
  40119, 40150,
  40150, 40181,
  40181, 40209,
  40209, 40240,
  40240, 40270,
  40270, 40301,
  40301, 40331,
  40331, 40362,
  40362, 40393,
  40393, 40423,
  40423, 40454,
  40454, 40484,
  40484, 40515,
  40515, 40546,
  40546, 40574,
  40574, 40605,
  40605, 40635,
  40635, 40666,
  40666, 40696,
  40696, 40727,
  40727, 40758,
  40758, 40788,
  40788, 40819,
  40819, 40849,
  40849, 40880,
  40880, 40911,
  40911, 40939,
  40939, 40970,
  40970, 41000,
  41000, 41031,
  41031, 41061,
  41061, 41092,
  41092, 41123,
  41123, 41153,
  41153, 41184,
  41184, 41214,
  41214, 41245,
  41245, 41276,
  41276, 41304,
  41304, 41335,
  41335, 41365,
  41365, 41396,
  41396, 41426,
  41426, 41457,
  41457, 41488,
  41488, 41518,
  41518, 41549,
  41549, 41579,
  41579, 41610,
  41610, 41641,
  41641, 41669,
  41669, 41700,
  41700, 41730,
  41730, 41761,
  41761, 41791,
  41791, 41822,
  41822, 41853,
  41853, 41883,
  41883, 41914,
  41914, 41944,
  41944, 41975,
  41975, 42006,
  42006, 42034,
  42034, 42065,
  42065, 42095,
  42095, 42126,
  42126, 42156,
  42156, 42187,
  42187, 42218,
  42218, 42248,
  42248, 42279,
  42279, 42309,
  42309, 42340,
  42340, 42371,
  42371, 42399,
  42399, 42430,
  42430, 42460,
  42460, 42491,
  42491, 42521,
  42521, 42552,
  42552, 42583,
  42583, 42613,
  42613, 42644,
  42644, 42674,
  42674, 42705,
  42705, 42736,
  42736, 42764,
  42764, 42795,
  42795, 42825,
  42825, 42856,
  42856, 42886,
  42886, 42917,
  42917, 42948,
  42948, 42978,
  42978, 43009,
  43009, 43039,
  43039, 43070,
  43070, 43101,
  43101, 43129,
  43129, 43160,
  43160, 43190,
  43190, 43221,
  43221, 43251,
  43251, 43282,
  43282, 43313,
  43313, 43343,
  43343, 43374,
  43374, 43404,
  43404, 43435,
  43435, 43466,
  43466, 43494,
  43494, 43525,
  43525, 43555,
  43555, 43586,
  43586, 43616,
  43616, 43647,
  43647, 43678,
  43678, 43708,
  43708, 43739,
  43739, 43769,
  43769, 43800,
  43800, 43831,
  43831, 43859,
  43859, 43890,
  43890, 43920,
  43920, 43951,
  43951, 43981,
  43981, 44012,
  44012, 44043,
  44043, 44073,
  44073, 44104,
  44104, 44134,
  44134, 44165,
  44165, 44196,
  44196, 44224,
  44224, 44255,
  44255, 44285,
  44285, 44316,
  44316, 44346,
  44346, 44377,
  44377, 44408,
  44408, 44438,
  44438, 44469,
  44469, 44499,
  44499, 44530,
  44530, 44561,
  44561, 44589,
  44589, 44620,
  44620, 44650,
  44650, 44681,
  44681, 44711,
  44711, 44742,
  44742, 44773,
  44773, 44803,
  44803, 44834,
  44834, 44864,
  44864, 44895,
  44895, 44926,
  44926, 44954,
  44954, 44985,
  44985, 45015,
  45015, 45046,
  45046, 45076,
  45076, 45107,
  45107, 45138,
  45138, 45168,
  45168, 45199,
  45199, 45229,
  45229, 45260,
  45260, 45291,
  45291, 45319,
  45319, 45350,
  45350, 45380,
  45380, 45411,
  45411, 45441,
  45441, 45472,
  45472, 45503,
  45503, 45533,
  45533, 45564,
  45564, 45594,
  45594, 45625,
  45625, 45656,
  45656, 45684,
  45684, 45715,
  45715, 45745,
  45745, 45776,
  45776, 45806,
  45806, 45837,
  45837, 45868,
  45868, 45898,
  45898, 45929,
  45929, 45959,
  45959, 45990,
  45990, 46021,
  46021, 46049,
  46049, 46080,
  46080, 46110,
  46110, 46141,
  46141, 46171,
  46171, 46202,
  46202, 46233,
  46233, 46263,
  46263, 46294,
  46294, 46324,
  46324, 46355,
  46355, 46386,
  46386, 46414,
  46414, 46445,
  46445, 46475,
  46475, 46506,
  46506, 46536,
  46536, 46567,
  46567, 46598,
  46598, 46628,
  46628, 46659,
  46659, 46689,
  46689, 46720,
  46720, 46751,
  46751, 46779,
  46779, 46810,
  46810, 46840,
  46840, 46871,
  46871, 46901,
  46901, 46932,
  46932, 46963,
  46963, 46993,
  46993, 47024,
  47024, 47054,
  47054, 47085,
  47085, 47116,
  47116, 47144,
  47144, 47175,
  47175, 47205,
  47205, 47236,
  47236, 47266,
  47266, 47297,
  47297, 47328,
  47328, 47358,
  47358, 47389,
  47389, 47419,
  47419, 47450,
  47450, 47481,
  47481, 47509,
  47509, 47540,
  47540, 47570,
  47570, 47601,
  47601, 47631,
  47631, 47662,
  47662, 47693,
  47693, 47723,
  47723, 47754,
  47754, 47784,
  47784, 47815,
  47815, 47846,
  47846, 47874,
  47874, 47905,
  47905, 47935,
  47935, 47966,
  47966, 47996,
  47996, 48027,
  48027, 48058,
  48058, 48088,
  48088, 48119,
  48119, 48149,
  48149, 48180,
  48180, 48211,
  48211, 48239,
  48239, 48270,
  48270, 48300,
  48300, 48331,
  48331, 48361,
  48361, 48392,
  48392, 48423,
  48423, 48453,
  48453, 48484,
  48484, 48514,
  48514, 48545,
  48545, 48576,
  48576, 48604,
  48604, 48635,
  48635, 48665,
  48665, 48696,
  48696, 48726,
  48726, 48757,
  48757, 48788,
  48788, 48818,
  48818, 48849,
  48849, 48879,
  48879, 48910,
  48910, 48941,
  48941, 48969,
  48969, 49000,
  49000, 49030,
  49030, 49061,
  49061, 49091,
  49091, 49122,
  49122, 49153,
  49153, 49183,
  49183, 49214,
  49214, 49244,
  49244, 49275,
  49275, 49306,
  49306, 49334,
  49334, 49365,
  49365, 49395,
  49395, 49426,
  49426, 49456,
  49456, 49487,
  49487, 49518,
  49518, 49548,
  49548, 49579,
  49579, 49609,
  49609, 49640,
  49640, 49671,
  49671, 49699,
  49699, 49730,
  49730, 49760,
  49760, 49791,
  49791, 49821,
  49821, 49852,
  49852, 49883,
  49883, 49913,
  49913, 49944,
  49944, 49974,
  49974, 50005,
  50005, 50036,
  50036, 50064,
  50064, 50095,
  50095, 50125,
  50125, 50156,
  50156, 50186,
  50186, 50217,
  50217, 50248,
  50248, 50278,
  50278, 50309,
  50309, 50339,
  50339, 50370,
  50370, 50401,
  50401, 50429,
  50429, 50460,
  50460, 50490,
  50490, 50521,
  50521, 50551,
  50551, 50582,
  50582, 50613,
  50613, 50643,
  50643, 50674,
  50674, 50704,
  50704, 50735,
  50735, 50766,
  50766, 50794,
  50794, 50825,
  50825, 50855,
  50855, 50886,
  50886, 50916,
  50916, 50947,
  50947, 50978,
  50978, 51008,
  51008, 51039,
  51039, 51069,
  51069, 51100,
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;

 lat = _ ;

 lon = _ ;

 z = _ ;

 temperature =
  _, _,
  _, _,
  _, _,
  _, _ ;
}
