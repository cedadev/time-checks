netcdf test_mon_360_day {
dimensions:
	time = UNLIMITED ;
	lat = 2 ;
	lon = 2 ;
    bnds = 2 ;
variables:
	double time(time) ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1859-12-01" ;
		time:calendar = "360_day" ;
		time:axis = "T" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
	double time_bnds(time, bnds) ;
	float lat ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "Latitude" ;
	float lon ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "Longitude" ;
	float z ;
		z:standard_name = "depth" ;
		z:positive = "down" ;
		z:units = "m" ;
		z:long_name = "Depth below surface" ;
	float temperature(time, lat, lon) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "deg_C" ;
		temperature:long_name = "Seawater Temperature" ;
		temperature:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:variable_id = "temp-max" ;
		:scenario = "sres-a1b" ;
		:dataset_id = "ukcp18-land-prob-25km" ;
		:prob_type = "sample" ;
		:frequency = "mon" ;
data:

 time = 18015, 18045, 18075, 18105, 18135, 18165, 18195, 18225, 18255, 18285,
    18315, 18345, 18375, 18405, 18435, 18465, 18495, 18525, 18555, 18585,
    18615, 18645, 18675, 18705, 18735, 18765, 18795, 18825, 18855, 18885,
    18915, 18945, 18975, 19005, 19035, 19065, 19095, 19125, 19155, 19185,
    19215, 19245, 19275, 19305, 19335, 19365, 19395, 19425, 19455, 19485,
    19515, 19545, 19575, 19605, 19635, 19665, 19695, 19725, 19755, 19785,
    19815, 19845, 19875, 19905, 19935, 19965, 19995, 20025, 20055, 20085,
    20115, 20145, 20175, 20205, 20235, 20265, 20295, 20325, 20355, 20385,
    20415, 20445, 20475, 20505, 20535, 20565, 20595, 20625, 20655, 20685,
    20715, 20745, 20775, 20805, 20835, 20865, 20895, 20925, 20955, 20985,
    21015, 21045, 21075, 21105, 21135, 21165, 21195, 21225, 21255, 21285,
    21315, 21345, 21375, 21405, 21435, 21465, 21495, 21525, 21555, 21585,
    21615, 21645, 21675, 21705, 21735, 21765, 21795, 21825, 21855, 21885,
    21915, 21945, 21975, 22005, 22035, 22065, 22095, 22125, 22155, 22185,
    22215, 22245, 22275, 22305, 22335, 22365, 22395, 22425, 22455, 22485,
    22515, 22545, 22575, 22605, 22635, 22665, 22695, 22725, 22755, 22785,
    22815, 22845, 22875, 22905, 22935, 22965, 22995, 23025, 23055, 23085,
    23115, 23145, 23175, 23205, 23235, 23265, 23295, 23325, 23355, 23385,
    23415, 23445, 23475, 23505, 23535, 23565, 23595, 23625, 23655, 23685,
    23715, 23745, 23775, 23805, 23835, 23865, 23895, 23925, 23955, 23985,
    24015, 24045, 24075, 24105, 24135, 24165, 24195, 24225, 24255, 24285,
    24315, 24345, 24375, 24405, 24435, 24465, 24495, 24525, 24555, 24585,
    24615, 24645, 24675, 24705, 24735, 24765, 24795, 24825, 24855, 24885,
    24915, 24945, 24975, 25005, 25035, 25065, 25095, 25125, 25155, 25185,
    25215, 25245, 25275, 25305, 25335, 25365, 25395, 25425, 25455, 25485,
    25515, 25545, 25575, 25605, 25635, 25665, 25695, 25725, 25755, 25785,
    25815, 25845, 25875, 25905, 25935, 25965, 25995, 26025, 26055, 26085,
    26115, 26145, 26175, 26205, 26235, 26265, 26295, 26325, 26355, 26385,
    26415, 26445, 26475, 26505, 26535, 26565, 26595, 26625, 26655, 26685,
    26715, 26745, 26775, 26805, 26835, 26865, 26895, 26925, 26955, 26985 ;

 time_bnds =
  18000, 18030,
  18030, 18060,
  18060, 18090,
  18090, 18120,
  18120, 18150,
  18150, 18180,
  18180, 18210,
  18210, 18240,
  18240, 18270,
  18270, 18300,
  18300, 18330,
  18330, 18360,
  18360, 18390,
  18390, 18420,
  18420, 18450,
  18450, 18480,
  18480, 18510,
  18510, 18540,
  18540, 18570,
  18570, 18600,
  18600, 18630,
  18630, 18660,
  18660, 18690,
  18690, 18720,
  18720, 18750,
  18750, 18780,
  18780, 18810,
  18810, 18840,
  18840, 18870,
  18870, 18900,
  18900, 18930,
  18930, 18960,
  18960, 18990,
  18990, 19020,
  19020, 19050,
  19050, 19080,
  19080, 19110,
  19110, 19140,
  19140, 19170,
  19170, 19200,
  19200, 19230,
  19230, 19260,
  19260, 19290,
  19290, 19320,
  19320, 19350,
  19350, 19380,
  19380, 19410,
  19410, 19440,
  19440, 19470,
  19470, 19500,
  19500, 19530,
  19530, 19560,
  19560, 19590,
  19590, 19620,
  19620, 19650,
  19650, 19680,
  19680, 19710,
  19710, 19740,
  19740, 19770,
  19770, 19800,
  19800, 19830,
  19830, 19860,
  19860, 19890,
  19890, 19920,
  19920, 19950,
  19950, 19980,
  19980, 20010,
  20010, 20040,
  20040, 20070,
  20070, 20100,
  20100, 20130,
  20130, 20160,
  20160, 20190,
  20190, 20220,
  20220, 20250,
  20250, 20280,
  20280, 20310,
  20310, 20340,
  20340, 20370,
  20370, 20400,
  20400, 20430,
  20430, 20460,
  20460, 20490,
  20490, 20520,
  20520, 20550,
  20550, 20580,
  20580, 20610,
  20610, 20640,
  20640, 20670,
  20670, 20700,
  20700, 20730,
  20730, 20760,
  20760, 20790,
  20790, 20820,
  20820, 20850,
  20850, 20880,
  20880, 20910,
  20910, 20940,
  20940, 20970,
  20970, 21000,
  21000, 21030,
  21030, 21060,
  21060, 21090,
  21090, 21120,
  21120, 21150,
  21150, 21180,
  21180, 21210,
  21210, 21240,
  21240, 21270,
  21270, 21300,
  21300, 21330,
  21330, 21360,
  21360, 21390,
  21390, 21420,
  21420, 21450,
  21450, 21480,
  21480, 21510,
  21510, 21540,
  21540, 21570,
  21570, 21600,
  21600, 21630,
  21630, 21660,
  21660, 21690,
  21690, 21720,
  21720, 21750,
  21750, 21780,
  21780, 21810,
  21810, 21840,
  21840, 21870,
  21870, 21900,
  21900, 21930,
  21930, 21960,
  21960, 21990,
  21990, 22020,
  22020, 22050,
  22050, 22080,
  22080, 22110,
  22110, 22140,
  22140, 22170,
  22170, 22200,
  22200, 22230,
  22230, 22260,
  22260, 22290,
  22290, 22320,
  22320, 22350,
  22350, 22380,
  22380, 22410,
  22410, 22440,
  22440, 22470,
  22470, 22500,
  22500, 22530,
  22530, 22560,
  22560, 22590,
  22590, 22620,
  22620, 22650,
  22650, 22680,
  22680, 22710,
  22710, 22740,
  22740, 22770,
  22770, 22800,
  22800, 22830,
  22830, 22860,
  22860, 22890,
  22890, 22920,
  22920, 22950,
  22950, 22980,
  22980, 23010,
  23010, 23040,
  23040, 23070,
  23070, 23100,
  23100, 23130,
  23130, 23160,
  23160, 23190,
  23190, 23220,
  23220, 23250,
  23250, 23280,
  23280, 23310,
  23310, 23340,
  23340, 23370,
  23370, 23400,
  23400, 23430,
  23430, 23460,
  23460, 23490,
  23490, 23520,
  23520, 23550,
  23550, 23580,
  23580, 23610,
  23610, 23640,
  23640, 23670,
  23670, 23700,
  23700, 23730,
  23730, 23760,
  23760, 23790,
  23790, 23820,
  23820, 23850,
  23850, 23880,
  23880, 23910,
  23910, 23940,
  23940, 23970,
  23970, 24000,
  24000, 24030,
  24030, 24060,
  24060, 24090,
  24090, 24120,
  24120, 24150,
  24150, 24180,
  24180, 24210,
  24210, 24240,
  24240, 24270,
  24270, 24300,
  24300, 24330,
  24330, 24360,
  24360, 24390,
  24390, 24420,
  24420, 24450,
  24450, 24480,
  24480, 24510,
  24510, 24540,
  24540, 24570,
  24570, 24600,
  24600, 24630,
  24630, 24660,
  24660, 24690,
  24690, 24720,
  24720, 24750,
  24750, 24780,
  24780, 24810,
  24810, 24840,
  24840, 24870,
  24870, 24900,
  24900, 24930,
  24930, 24960,
  24960, 24990,
  24990, 25020,
  25020, 25050,
  25050, 25080,
  25080, 25110,
  25110, 25140,
  25140, 25170,
  25170, 25200,
  25200, 25230,
  25230, 25260,
  25260, 25290,
  25290, 25320,
  25320, 25350,
  25350, 25380,
  25380, 25410,
  25410, 25440,
  25440, 25470,
  25470, 25500,
  25500, 25530,
  25530, 25560,
  25560, 25590,
  25590, 25620,
  25620, 25650,
  25650, 25680,
  25680, 25710,
  25710, 25740,
  25740, 25770,
  25770, 25800,
  25800, 25830,
  25830, 25860,
  25860, 25890,
  25890, 25920,
  25920, 25950,
  25950, 25980,
  25980, 26010,
  26010, 26040,
  26040, 26070,
  26070, 26100,
  26100, 26130,
  26130, 26160,
  26160, 26190,
  26190, 26220,
  26220, 26250,
  26250, 26280,
  26280, 26310,
  26310, 26340,
  26340, 26370,
  26370, 26400,
  26400, 26430,
  26430, 26460,
  26460, 26490,
  26490, 26520,
  26520, 26550,
  26550, 26580,
  26580, 26610,
  26610, 26640,
  26640, 26670,
  26670, 26700,
  26700, 26730,
  26730, 26760,
  26760, 26790,
  26790, 26820,
  26820, 26850,
  26850, 26880,
  26880, 26910,
  26910, 26940,
  26940, 26970,
  26970, 27000 ;

 lat = _ ;

 lon = _ ;

 z = _ ;

 temperature =
  _, _,
  _, _,
  _, _,
  _, _ ;
}
