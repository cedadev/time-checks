netcdf test_mon_gregorian {
dimensions:
	time = UNLIMITED ;
	lat = 2 ;
	lon = 2 ;
    bnds = 2 ;
variables:
	double time(time) ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1850-1-1" ;
		time:calendar = "gregorian" ;
		time:axis = "T" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
	double time_bnds(time, bnds) ;
	float lat ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "Latitude" ;
	float lon ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "Longitude" ;
	float z ;
		z:standard_name = "depth" ;
		z:positive = "down" ;
		z:units = "m" ;
		z:long_name = "Depth below surface" ;
	float temperature(time, lat, lon) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "deg_C" ;
		temperature:long_name = "Seawater Temperature" ;
		temperature:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:variable_id = "temp-max" ;
		:scenario = "sres-a1b" ;
		:dataset_id = "ukcp18-land-prob-25km" ;
		:prob_type = "sample" ;
		:frequency = "mon" ;
data:

 time = 18277.5, 18307, 18336.5, 18367, 18397.5, 18428, 18458.5, 18489.5,
    18520, 18550.5, 18581, 18611.5, 18642.5, 18672, 18701.5, 18732, 18762.5,
    18793, 18823.5, 18854.5, 18885, 18915.5, 18946, 18976.5, 19007.5, 19037,
    19066.5, 19097, 19127.5, 19158, 19188.5, 19219.5, 19250, 19280.5, 19311,
    19341.5, 19372.5, 19402, 19431.5, 19462, 19492.5, 19523, 19553.5,
    19584.5, 19615, 19645.5, 19676, 19706.5, 19737.5, 19767.5, 19797.5,
    19828, 19858.5, 19889, 19919.5, 19950.5, 19981, 20011.5, 20042, 20072.5,
    20103.5, 20133, 20162.5, 20193, 20223.5, 20254, 20284.5, 20315.5, 20346,
    20376.5, 20407, 20437.5, 20468.5, 20498, 20527.5, 20558, 20588.5, 20619,
    20649.5, 20680.5, 20711, 20741.5, 20772, 20802.5, 20833.5, 20863,
    20892.5, 20923, 20953.5, 20984, 21014.5, 21045.5, 21076, 21106.5, 21137,
    21167.5, 21198.5, 21228.5, 21258.5, 21289, 21319.5, 21350, 21380.5,
    21411.5, 21442, 21472.5, 21503, 21533.5, 21564.5, 21594, 21623.5, 21654,
    21684.5, 21715, 21745.5, 21776.5, 21807, 21837.5, 21868, 21898.5,
    21929.5, 21959, 21988.5, 22019, 22049.5, 22080, 22110.5, 22141.5, 22172,
    22202.5, 22233, 22263.5, 22294.5, 22324, 22353.5, 22384, 22414.5, 22445,
    22475.5, 22506.5, 22537, 22567.5, 22598, 22628.5, 22659.5, 22689.5,
    22719.5, 22750, 22780.5, 22811, 22841.5, 22872.5, 22903, 22933.5, 22964,
    22994.5, 23025.5, 23055, 23084.5, 23115, 23145.5, 23176, 23206.5,
    23237.5, 23268, 23298.5, 23329, 23359.5, 23390.5, 23420, 23449.5, 23480,
    23510.5, 23541, 23571.5, 23602.5, 23633, 23663.5, 23694, 23724.5,
    23755.5, 23785, 23814.5, 23845, 23875.5, 23906, 23936.5, 23967.5, 23998,
    24028.5, 24059, 24089.5, 24120.5, 24150.5, 24180.5, 24211, 24241.5,
    24272, 24302.5, 24333.5, 24364, 24394.5, 24425, 24455.5, 24486.5, 24516,
    24545.5, 24576, 24606.5, 24637, 24667.5, 24698.5, 24729, 24759.5, 24790,
    24820.5, 24851.5, 24881, 24910.5, 24941, 24971.5, 25002, 25032.5,
    25063.5, 25094, 25124.5, 25155, 25185.5, 25216.5, 25246, 25275.5, 25306,
    25336.5, 25367, 25397.5, 25428.5, 25459, 25489.5, 25520, 25550.5,
    25581.5, 25611.5, 25641.5, 25672, 25702.5, 25733, 25763.5, 25794.5,
    25825, 25855.5, 25886, 25916.5, 25947.5, 25977, 26006.5, 26037, 26067.5,
    26098, 26128.5, 26159.5, 26190, 26220.5, 26251, 26281.5, 26312.5, 26342,
    26371.5, 26402, 26432.5, 26463, 26493.5, 26524.5, 26555, 26585.5, 26616,
    26646.5, 26677.5, 26707, 26736.5, 26767, 26797.5, 26828, 26858.5,
    26889.5, 26920, 26950.5, 26981, 27011.5, 27042.5, 27072.5, 27102.5,
    27133, 27163.5, 27194, 27224.5, 27255.5, 27286, 27316.5, 27347, 27377.5,
    27408.5, 27438, 27467.5, 27498, 27528.5, 27559, 27589.5, 27620.5, 27651,
    27681.5, 27712, 27742.5, 27773.5, 27803, 27832.5, 27863, 27893.5, 27924,
    27954.5, 27985.5, 28016, 28046.5, 28077, 28107.5, 28138.5, 28168,
    28197.5, 28228, 28258.5, 28289, 28319.5, 28350.5, 28381, 28411.5, 28442,
    28472.5, 28503.5, 28533.5, 28563.5, 28594, 28624.5, 28655, 28685.5,
    28716.5, 28747, 28777.5, 28808, 28838.5, 28869.5, 28899, 28928.5, 28959,
    28989.5, 29020, 29050.5, 29081.5, 29112, 29142.5, 29173, 29203.5,
    29234.5, 29264, 29293.5, 29324, 29354.5, 29385, 29415.5, 29446.5, 29477,
    29507.5, 29538, 29568.5, 29599.5, 29629, 29658.5, 29689, 29719.5, 29750,
    29780.5, 29811.5, 29842, 29872.5, 29903, 29933.5, 29964.5, 29994.5,
    30024.5, 30055, 30085.5, 30116, 30146.5, 30177.5, 30208, 30238.5, 30269,
    30299.5, 30330.5, 30360, 30389.5, 30420, 30450.5, 30481, 30511.5,
    30542.5, 30573, 30603.5, 30634, 30664.5, 30695.5, 30725, 30754.5, 30785,
    30815.5, 30846, 30876.5, 30907.5, 30938, 30968.5, 30999, 31029.5,
    31060.5, 31090, 31119.5, 31150, 31180.5, 31211, 31241.5, 31272.5, 31303,
    31333.5, 31364, 31394.5, 31425.5, 31455.5, 31485.5, 31516, 31546.5,
    31577, 31607.5, 31638.5, 31669, 31699.5, 31730, 31760.5, 31791.5, 31821,
    31850.5, 31881, 31911.5, 31942, 31972.5, 32003.5, 32034, 32064.5, 32095,
    32125.5, 32156.5, 32186, 32215.5, 32246, 32276.5, 32307, 32337.5,
    32368.5, 32399, 32429.5, 32460, 32490.5, 32521.5, 32551, 32580.5, 32611,
    32641.5, 32672, 32702.5, 32733.5, 32764, 32794.5, 32825, 32855.5,
    32886.5, 32916.5, 32946.5, 32977, 33007.5, 33038, 33068.5, 33099.5,
    33130, 33160.5, 33191, 33221.5, 33252.5, 33282, 33311.5, 33342, 33372.5,
    33403, 33433.5, 33464.5, 33495, 33525.5, 33556, 33586.5, 33617.5, 33647,
    33676.5, 33707, 33737.5, 33768, 33798.5, 33829.5, 33860, 33890.5, 33921,
    33951.5, 33982.5, 34012, 34041.5, 34072, 34102.5, 34133, 34163.5,
    34194.5, 34225, 34255.5, 34286, 34316.5, 34347.5, 34377.5, 34407.5,
    34438, 34468.5, 34499, 34529.5, 34560.5, 34591, 34621.5, 34652, 34682.5,
    34713.5, 34743, 34772.5, 34803, 34833.5, 34864, 34894.5, 34925.5, 34956,
    34986.5, 35017, 35047.5, 35078.5, 35108, 35137.5, 35168, 35198.5, 35229,
    35259.5, 35290.5, 35321, 35351.5, 35382, 35412.5, 35443.5, 35473,
    35502.5, 35533, 35563.5, 35594, 35624.5, 35655.5, 35686, 35716.5, 35747,
    35777.5, 35808.5, 35838.5, 35868.5, 35899, 35929.5, 35960, 35990.5,
    36021.5, 36052, 36082.5, 36113, 36143.5, 36174.5, 36204, 36233.5, 36264,
    36294.5, 36325, 36355.5, 36386.5, 36417, 36447.5, 36478, 36508.5 ;

 time_bnds =
  18262, 18293,
  18293, 18321,
  18321, 18352,
  18352, 18382,
  18382, 18413,
  18413, 18443,
  18443, 18474,
  18474, 18505,
  18505, 18535,
  18535, 18566,
  18566, 18596,
  18596, 18627,
  18627, 18658,
  18658, 18686,
  18686, 18717,
  18717, 18747,
  18747, 18778,
  18778, 18808,
  18808, 18839,
  18839, 18870,
  18870, 18900,
  18900, 18931,
  18931, 18961,
  18961, 18992,
  18992, 19023,
  19023, 19051,
  19051, 19082,
  19082, 19112,
  19112, 19143,
  19143, 19173,
  19173, 19204,
  19204, 19235,
  19235, 19265,
  19265, 19296,
  19296, 19326,
  19326, 19357,
  19357, 19388,
  19388, 19416,
  19416, 19447,
  19447, 19477,
  19477, 19508,
  19508, 19538,
  19538, 19569,
  19569, 19600,
  19600, 19630,
  19630, 19661,
  19661, 19691,
  19691, 19722,
  19722, 19753,
  19753, 19782,
  19782, 19813,
  19813, 19843,
  19843, 19874,
  19874, 19904,
  19904, 19935,
  19935, 19966,
  19966, 19996,
  19996, 20027,
  20027, 20057,
  20057, 20088,
  20088, 20119,
  20119, 20147,
  20147, 20178,
  20178, 20208,
  20208, 20239,
  20239, 20269,
  20269, 20300,
  20300, 20331,
  20331, 20361,
  20361, 20392,
  20392, 20422,
  20422, 20453,
  20453, 20484,
  20484, 20512,
  20512, 20543,
  20543, 20573,
  20573, 20604,
  20604, 20634,
  20634, 20665,
  20665, 20696,
  20696, 20726,
  20726, 20757,
  20757, 20787,
  20787, 20818,
  20818, 20849,
  20849, 20877,
  20877, 20908,
  20908, 20938,
  20938, 20969,
  20969, 20999,
  20999, 21030,
  21030, 21061,
  21061, 21091,
  21091, 21122,
  21122, 21152,
  21152, 21183,
  21183, 21214,
  21214, 21243,
  21243, 21274,
  21274, 21304,
  21304, 21335,
  21335, 21365,
  21365, 21396,
  21396, 21427,
  21427, 21457,
  21457, 21488,
  21488, 21518,
  21518, 21549,
  21549, 21580,
  21580, 21608,
  21608, 21639,
  21639, 21669,
  21669, 21700,
  21700, 21730,
  21730, 21761,
  21761, 21792,
  21792, 21822,
  21822, 21853,
  21853, 21883,
  21883, 21914,
  21914, 21945,
  21945, 21973,
  21973, 22004,
  22004, 22034,
  22034, 22065,
  22065, 22095,
  22095, 22126,
  22126, 22157,
  22157, 22187,
  22187, 22218,
  22218, 22248,
  22248, 22279,
  22279, 22310,
  22310, 22338,
  22338, 22369,
  22369, 22399,
  22399, 22430,
  22430, 22460,
  22460, 22491,
  22491, 22522,
  22522, 22552,
  22552, 22583,
  22583, 22613,
  22613, 22644,
  22644, 22675,
  22675, 22704,
  22704, 22735,
  22735, 22765,
  22765, 22796,
  22796, 22826,
  22826, 22857,
  22857, 22888,
  22888, 22918,
  22918, 22949,
  22949, 22979,
  22979, 23010,
  23010, 23041,
  23041, 23069,
  23069, 23100,
  23100, 23130,
  23130, 23161,
  23161, 23191,
  23191, 23222,
  23222, 23253,
  23253, 23283,
  23283, 23314,
  23314, 23344,
  23344, 23375,
  23375, 23406,
  23406, 23434,
  23434, 23465,
  23465, 23495,
  23495, 23526,
  23526, 23556,
  23556, 23587,
  23587, 23618,
  23618, 23648,
  23648, 23679,
  23679, 23709,
  23709, 23740,
  23740, 23771,
  23771, 23799,
  23799, 23830,
  23830, 23860,
  23860, 23891,
  23891, 23921,
  23921, 23952,
  23952, 23983,
  23983, 24013,
  24013, 24044,
  24044, 24074,
  24074, 24105,
  24105, 24136,
  24136, 24165,
  24165, 24196,
  24196, 24226,
  24226, 24257,
  24257, 24287,
  24287, 24318,
  24318, 24349,
  24349, 24379,
  24379, 24410,
  24410, 24440,
  24440, 24471,
  24471, 24502,
  24502, 24530,
  24530, 24561,
  24561, 24591,
  24591, 24622,
  24622, 24652,
  24652, 24683,
  24683, 24714,
  24714, 24744,
  24744, 24775,
  24775, 24805,
  24805, 24836,
  24836, 24867,
  24867, 24895,
  24895, 24926,
  24926, 24956,
  24956, 24987,
  24987, 25017,
  25017, 25048,
  25048, 25079,
  25079, 25109,
  25109, 25140,
  25140, 25170,
  25170, 25201,
  25201, 25232,
  25232, 25260,
  25260, 25291,
  25291, 25321,
  25321, 25352,
  25352, 25382,
  25382, 25413,
  25413, 25444,
  25444, 25474,
  25474, 25505,
  25505, 25535,
  25535, 25566,
  25566, 25597,
  25597, 25626,
  25626, 25657,
  25657, 25687,
  25687, 25718,
  25718, 25748,
  25748, 25779,
  25779, 25810,
  25810, 25840,
  25840, 25871,
  25871, 25901,
  25901, 25932,
  25932, 25963,
  25963, 25991,
  25991, 26022,
  26022, 26052,
  26052, 26083,
  26083, 26113,
  26113, 26144,
  26144, 26175,
  26175, 26205,
  26205, 26236,
  26236, 26266,
  26266, 26297,
  26297, 26328,
  26328, 26356,
  26356, 26387,
  26387, 26417,
  26417, 26448,
  26448, 26478,
  26478, 26509,
  26509, 26540,
  26540, 26570,
  26570, 26601,
  26601, 26631,
  26631, 26662,
  26662, 26693,
  26693, 26721,
  26721, 26752,
  26752, 26782,
  26782, 26813,
  26813, 26843,
  26843, 26874,
  26874, 26905,
  26905, 26935,
  26935, 26966,
  26966, 26996,
  26996, 27027,
  27027, 27058,
  27058, 27087,
  27087, 27118,
  27118, 27148,
  27148, 27179,
  27179, 27209,
  27209, 27240,
  27240, 27271,
  27271, 27301,
  27301, 27332,
  27332, 27362,
  27362, 27393,
  27393, 27424,
  27424, 27452,
  27452, 27483,
  27483, 27513,
  27513, 27544,
  27544, 27574,
  27574, 27605,
  27605, 27636,
  27636, 27666,
  27666, 27697,
  27697, 27727,
  27727, 27758,
  27758, 27789,
  27789, 27817,
  27817, 27848,
  27848, 27878,
  27878, 27909,
  27909, 27939,
  27939, 27970,
  27970, 28001,
  28001, 28031,
  28031, 28062,
  28062, 28092,
  28092, 28123,
  28123, 28154,
  28154, 28182,
  28182, 28213,
  28213, 28243,
  28243, 28274,
  28274, 28304,
  28304, 28335,
  28335, 28366,
  28366, 28396,
  28396, 28427,
  28427, 28457,
  28457, 28488,
  28488, 28519,
  28519, 28548,
  28548, 28579,
  28579, 28609,
  28609, 28640,
  28640, 28670,
  28670, 28701,
  28701, 28732,
  28732, 28762,
  28762, 28793,
  28793, 28823,
  28823, 28854,
  28854, 28885,
  28885, 28913,
  28913, 28944,
  28944, 28974,
  28974, 29005,
  29005, 29035,
  29035, 29066,
  29066, 29097,
  29097, 29127,
  29127, 29158,
  29158, 29188,
  29188, 29219,
  29219, 29250,
  29250, 29278,
  29278, 29309,
  29309, 29339,
  29339, 29370,
  29370, 29400,
  29400, 29431,
  29431, 29462,
  29462, 29492,
  29492, 29523,
  29523, 29553,
  29553, 29584,
  29584, 29615,
  29615, 29643,
  29643, 29674,
  29674, 29704,
  29704, 29735,
  29735, 29765,
  29765, 29796,
  29796, 29827,
  29827, 29857,
  29857, 29888,
  29888, 29918,
  29918, 29949,
  29949, 29980,
  29980, 30009,
  30009, 30040,
  30040, 30070,
  30070, 30101,
  30101, 30131,
  30131, 30162,
  30162, 30193,
  30193, 30223,
  30223, 30254,
  30254, 30284,
  30284, 30315,
  30315, 30346,
  30346, 30374,
  30374, 30405,
  30405, 30435,
  30435, 30466,
  30466, 30496,
  30496, 30527,
  30527, 30558,
  30558, 30588,
  30588, 30619,
  30619, 30649,
  30649, 30680,
  30680, 30711,
  30711, 30739,
  30739, 30770,
  30770, 30800,
  30800, 30831,
  30831, 30861,
  30861, 30892,
  30892, 30923,
  30923, 30953,
  30953, 30984,
  30984, 31014,
  31014, 31045,
  31045, 31076,
  31076, 31104,
  31104, 31135,
  31135, 31165,
  31165, 31196,
  31196, 31226,
  31226, 31257,
  31257, 31288,
  31288, 31318,
  31318, 31349,
  31349, 31379,
  31379, 31410,
  31410, 31441,
  31441, 31470,
  31470, 31501,
  31501, 31531,
  31531, 31562,
  31562, 31592,
  31592, 31623,
  31623, 31654,
  31654, 31684,
  31684, 31715,
  31715, 31745,
  31745, 31776,
  31776, 31807,
  31807, 31835,
  31835, 31866,
  31866, 31896,
  31896, 31927,
  31927, 31957,
  31957, 31988,
  31988, 32019,
  32019, 32049,
  32049, 32080,
  32080, 32110,
  32110, 32141,
  32141, 32172,
  32172, 32200,
  32200, 32231,
  32231, 32261,
  32261, 32292,
  32292, 32322,
  32322, 32353,
  32353, 32384,
  32384, 32414,
  32414, 32445,
  32445, 32475,
  32475, 32506,
  32506, 32537,
  32537, 32565,
  32565, 32596,
  32596, 32626,
  32626, 32657,
  32657, 32687,
  32687, 32718,
  32718, 32749,
  32749, 32779,
  32779, 32810,
  32810, 32840,
  32840, 32871,
  32871, 32902,
  32902, 32931,
  32931, 32962,
  32962, 32992,
  32992, 33023,
  33023, 33053,
  33053, 33084,
  33084, 33115,
  33115, 33145,
  33145, 33176,
  33176, 33206,
  33206, 33237,
  33237, 33268,
  33268, 33296,
  33296, 33327,
  33327, 33357,
  33357, 33388,
  33388, 33418,
  33418, 33449,
  33449, 33480,
  33480, 33510,
  33510, 33541,
  33541, 33571,
  33571, 33602,
  33602, 33633,
  33633, 33661,
  33661, 33692,
  33692, 33722,
  33722, 33753,
  33753, 33783,
  33783, 33814,
  33814, 33845,
  33845, 33875,
  33875, 33906,
  33906, 33936,
  33936, 33967,
  33967, 33998,
  33998, 34026,
  34026, 34057,
  34057, 34087,
  34087, 34118,
  34118, 34148,
  34148, 34179,
  34179, 34210,
  34210, 34240,
  34240, 34271,
  34271, 34301,
  34301, 34332,
  34332, 34363,
  34363, 34392,
  34392, 34423,
  34423, 34453,
  34453, 34484,
  34484, 34514,
  34514, 34545,
  34545, 34576,
  34576, 34606,
  34606, 34637,
  34637, 34667,
  34667, 34698,
  34698, 34729,
  34729, 34757,
  34757, 34788,
  34788, 34818,
  34818, 34849,
  34849, 34879,
  34879, 34910,
  34910, 34941,
  34941, 34971,
  34971, 35002,
  35002, 35032,
  35032, 35063,
  35063, 35094,
  35094, 35122,
  35122, 35153,
  35153, 35183,
  35183, 35214,
  35214, 35244,
  35244, 35275,
  35275, 35306,
  35306, 35336,
  35336, 35367,
  35367, 35397,
  35397, 35428,
  35428, 35459,
  35459, 35487,
  35487, 35518,
  35518, 35548,
  35548, 35579,
  35579, 35609,
  35609, 35640,
  35640, 35671,
  35671, 35701,
  35701, 35732,
  35732, 35762,
  35762, 35793,
  35793, 35824,
  35824, 35853,
  35853, 35884,
  35884, 35914,
  35914, 35945,
  35945, 35975,
  35975, 36006,
  36006, 36037,
  36037, 36067,
  36067, 36098,
  36098, 36128,
  36128, 36159,
  36159, 36190,
  36190, 36218,
  36218, 36249,
  36249, 36279,
  36279, 36310,
  36310, 36340,
  36340, 36371,
  36371, 36402,
  36402, 36432,
  36432, 36463,
  36463, 36493,
  36493, 36524 ;

 lat = _ ;

 lon = _ ;

 z = _ ;

 temperature =
  _, _,
  _, _,
  _, _,
  _, _ ;
}
