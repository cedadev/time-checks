netcdf mrsos_day_HadGEM2-ES_historical_r1i1p1_19991201-20051130 {
dimensions:
	bnds = 2 ;
	lat = 2 ;
	lon = 2 ;
	time = UNLIMITED ; // (2160 currently)
variables:
	double depth ;
		depth:units = "m" ;
		depth:axis = "Z" ;
		depth:positive = "down" ;
		depth:long_name = "depth" ;
		depth:standard_name = "depth" ;
		depth:bounds = "depth_bnds" ;
	double depth_bnds(bnds) ;
	double lat(lat) ;
		lat:bounds = "lat_bnds" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:bounds = "lon_bnds" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
	double lon_bnds(lon, bnds) ;
	float mrsos(time, lat, lon) ;
		mrsos:standard_name = "moisture_content_of_soil_layer" ;
		mrsos:long_name = "Moisture in Upper 0.1 m of Soil Column" ;
		mrsos:comment = "Compute the mass of water in all phases in the upper 0.1 meters of soil." ;
		mrsos:units = "kg m-2" ;
		mrsos:original_name = "mo: m01s08i223" ;
		mrsos:cell_methods = "time: mean area: mean where land" ;
		mrsos:cell_measures = "area: areacella" ;
		mrsos:history = "2010-11-23T09:37:12Z altered by CMOR: Treated scalar dimension: \'depth\'. 2010-11-23T09:37:12Z altered by CMOR: replaced missing value flag (-1.07374e+09) with standard missing value (1e+20)." ;
		mrsos:coordinates = "depth" ;
		mrsos:missing_value = 1.e+20f ;
		mrsos:_FillValue = 1.e+20f ;
		mrsos:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_land_fx_HadGEM2-ES_historical_r0i0p0.nc areacella: areacella_fx_HadGEM2-ES_historical_r0i0p0.nc" ;
	double time(time) ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1859-12-01" ;
		time:calendar = "360_day" ;
		time:axis = "T" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:institution = "Met Office Hadley Centre, Fitzroy Road, Exeter, Devon, EX1 3PB, UK, (http://www.metoffice.gov.uk)" ;
		:institute_id = "MOHC" ;
		:experiment_id = "historical" ;
		:source = "HadGEM2-ES (2009) atmosphere: HadGAM2 (N96L38); ocean: HadGOM2 (lat: 1.0-0.3 lon: 1.0 L40); land-surface/vegetation: MOSES2 and TRIFFID; tropospheric chemistry: UKCA; ocean biogeochemistry: diat-HadOCC" ;
		:model_id = "HadGEM2-ES" ;
		:forcing = "GHG, SA, Oz, LU, Sl, Vl, BC, OC, (GHG = CO2, N2O, CH4, CFCs)" ;
		:parent_experiment_id = "piControl" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 0. ;
		:contact = "chris.d.jones@metoffice.gov.uk, michael.sanderson@metoffice.gov.uk" ;
		:history = "Wed Nov  1 09:35:58 2017: ncks -d lat,,,100 -d lon,,,100 -v mrsos /data/time-checks/mrsos_day_HadGEM2-ES_historical_r1i1p1_19991201-20051130.nc test_data/cmip5/mrsos_day_HadGEM2-ES_historical_r1i1p1_19991201-20051130.nc\n",
			"MOHC pp to CMOR/NetCDF convertor (version 1.5) 2010-11-23T09:37:09Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
		:references = "Bellouin N. et al, (2007) Improved representation of aerosols for HadGEM2. Meteorological Office Hadley Centre, Technical Note 73, March 2007; Collins W.J.  et al, (2008) Evaluation of the HadGEM2 model. Meteorological Office Hadley Centre, Technical Note 74,; Johns T.C. et al, (2006) The new Hadley Centre climate model HadGEM1: Evaluation of coupled simulations. Journal of Climate, American Meteorological Society, Vol. 19, No. 7, pages 1327-1353.; Martin G.M. et al, (2006) The physical properties of the atmosphere in the new Hadley Centre Global Environmental Model, HadGEM1 - Part 1: Model description and global climatology. Journal of Climate, American Meteorological Society, Vol. 19, No.7, pages 1274-1301.; Ringer M.A. et al, (2006) The physical properties of the atmosphere in the new Hadley Centre Global Environmental Model, HadGEM1 - Part 2: Aspects of variability and regional climate. Journal of Climate, American Meteorological Society, Vol. 19, No. 7, pages 1302-1326." ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "32d05752-0b67-44fd-b371-0c7fa22b400b" ;
		:mo_runid = "ajhoh" ;
		:product = "output" ;
		:experiment = "historical" ;
		:frequency = "day" ;
		:creation_date = "2010-11-23T11:30:25Z" ;
		:Conventions = "CF-1.4" ;
		:project_id = "CMIP5" ;
		:table_id = "Table day (12 November 2010) 53fa6f63b86081d1c644183416239052" ;
		:title = "HadGEM2-ES model output prepared for CMIP5 historical" ;
		:parent_experiment = "pre-industrial control" ;
		:modeling_realm = "land" ;
		:realization = 1 ;
		:cmor_version = "2.5.0" ;
		:NCO = "\"4.5.5\"" ;
data:

 depth = 0.05 ;

 depth_bnds = 0, 0.1 ;

 lat = -90, 35 ;

 lat_bnds =
  -90, -89.375,
  34.375, 35.625 ;

 lon = 0, 187.5 ;

 lon_bnds =
  -0.9375, 0.9375,
  186.5625, 188.4375 ;

 mrsos =
  0, 0,
  23.39478, _,
  0, 0,
  22.81311, _,
  0, 0,
  25.29138, _,
  0, 0,
  26.46545, _,
  0, 0,
  24.9751, _,
  0, 0,
  24.15149, _,
  0, 0,
  23.58478, _,
  0, 0,
  28.80652, _,
  0, 0,
  26.93085, _,
  0, 0,
  25.82062, _,
  0, 0,
  24.95587, _,
  0, 0,
  25.4447, _,
  0, 0,
  25.42444, _,
  0, 0,
  24.90204, _,
  0, 0,
  24.45428, _,
  0, 0,
  24.25116, _,
  0, 0,
  23.84918, _,
  0, 0,
  23.40961, _,
  0, 0,
  22.93689, _,
  0, 0,
  22.61426, _,
  0, 0,
  22.53839, _,
  0, 0,
  22.49371, _,
  0, 0,
  22.35339, _,
  0, 0,
  22.1095, _,
  0, 0,
  21.91895, _,
  0, 0,
  22.09985, _,
  0, 0,
  21.79254, _,
  0, 0,
  21.16132, _,
  0, 0,
  20.77167, _,
  0, 0,
  20.45752, _,
  0, 0,
  20.25012, _,
  0, 0,
  20.06952, _,
  0, 0,
  19.84674, _,
  0, 0,
  19.62909, _,
  0, 0,
  19.51959, _,
  0, 0,
  19.76819, _,
  0, 0,
  19.77246, _,
  0, 0,
  19.49023, _,
  0, 0,
  19.21216, _,
  0, 0,
  19.50543, _,
  0, 0,
  19.40448, _,
  0, 0,
  19.00671, _,
  0, 0,
  18.60071, _,
  0, 0,
  18.20355, _,
  0, 0,
  18.15967, _,
  0, 0,
  19.98169, _,
  0, 0,
  21.00519, _,
  0, 0,
  20.73407, _,
  0, 0,
  20.81476, _,
  0, 0,
  21.60034, _,
  0, 0,
  21.76392, _,
  0, 0,
  23.37872, _,
  0, 0,
  24.0708, _,
  0, 0,
  23.47028, _,
  0, 0,
  22.9071, _,
  0, 0,
  22.69751, _,
  0, 0,
  22.31543, _,
  0, 0,
  21.88556, _,
  0, 0,
  21.54651, _,
  0, 0,
  21.18658, _,
  0, 0,
  20.79407, _,
  0, 0,
  20.35516, _,
  0, 0,
  19.8183, _,
  0, 0,
  19.15912, _,
  0, 0,
  18.35156, _,
  0, 0,
  17.4295, _,
  0, 0,
  16.58356, _,
  0, 0,
  15.84558, _,
  0, 0,
  15.15997, _,
  0, 0,
  14.58154, _,
  0, 0,
  13.86798, _,
  0, 0,
  13.00671, _,
  0, 0,
  12.23956, _,
  0, 0,
  11.55408, _,
  0, 0,
  11.12909, _,
  0, 0,
  10.92719, _,
  0, 0,
  10.35382, _,
  0, 0,
  9.664551, _,
  0, 0,
  9.017029, _,
  0, 0,
  8.433472, _,
  0, 0,
  7.885071, _,
  0, 0,
  7.407898, _,
  0, 0,
  7.078613, _,
  0, 0,
  6.721375, _,
  0, 0,
  6.313599, _,
  0, 0,
  5.924194, _,
  0, 0,
  5.556702, _,
  0, 0,
  5.288147, _,
  0, 0,
  5.160828, _,
  0, 0,
  5.183533, _,
  0, 0,
  5.143005, _,
  0, 0,
  5.008545, _,
  0, 0,
  4.9729, _,
  0, 0,
  4.916504, _,
  0, 0,
  4.752441, _,
  0, 0,
  4.524414, _,
  0, 0,
  4.300598, _,
  0, 0,
  4.095581, _,
  0, 0,
  4.000183, _,
  0, 0,
  3.858093, _,
  0, 0,
  3.692444, _,
  0, 0,
  3.605835, _,
  0, 0,
  4.053528, _,
  0, 0,
  3.769287, _,
  0, 0,
  3.895203, _,
  0, 0,
  3.766357, _,
  0, 0,
  3.532104, _,
  0, 0,
  3.335815, _,
  0, 0,
  3.507507, _,
  0, 0,
  3.346069, _,
  0, 0,
  4.561829, _,
  0, 0,
  6.474121, _,
  0, 0,
  7.632446, _,
  0, 0,
  7.214539, _,
  0, 0,
  7.914429, _,
  0, 0,
  7.410095, _,
  0, 0,
  7.282837, _,
  0, 0,
  8.26001, _,
  0, 0,
  9.605225, _,
  0, 0,
  10.25378, _,
  0, 0,
  10.54626, _,
  0, 0,
  10.74115, _,
  0, 0,
  12.44592, _,
  0, 0,
  11.41138, _,
  0, 0,
  11.06396, _,
  0, 0,
  10.68579, _,
  0, 0,
  9.558105, _,
  0, 0,
  8.559143, _,
  0, 0,
  7.616516, _,
  0, 0,
  6.720825, _,
  0, 0,
  5.871521, _,
  0, 0,
  5.25354, _,
  0, 0,
  5.27594, _,
  0, 0,
  6.941467, _,
  0, 0,
  11.28961, _,
  0, 0,
  13.33606, _,
  0, 0,
  13.57861, _,
  0, 0,
  14.73938, _,
  0, 0,
  13.86218, _,
  0, 0,
  12.05707, _,
  0, 0,
  10.63947, _,
  0, 0,
  9.313232, _,
  0, 0,
  9.032959, _,
  0, 0,
  14.04578, _,
  0, 0,
  26.34375, _,
  0, 0,
  24.19623, _,
  0, 0,
  23.76685, _,
  0, 0,
  22.5528, _,
  0, 0,
  21.53784, _,
  0, 0,
  20.64111, _,
  0, 0,
  18.61603, _,
  0, 0,
  16.29352, _,
  0, 0,
  16.47473, _,
  0, 0,
  16.06543, _,
  0, 0,
  14.41016, _,
  0, 0,
  21.86597, _,
  0, 0,
  25.46692, _,
  0, 0,
  23.55371, _,
  0, 0,
  20.78845, _,
  0, 0,
  18.56177, _,
  0, 0,
  16.47455, _,
  0, 0,
  14.1131, _,
  0, 0,
  12.22742, _,
  0, 0,
  10.8147, _,
  0, 0,
  9.129883, _,
  0, 0,
  7.618896, _,
  0, 0,
  7.036499, _,
  0, 0,
  6.04126, _,
  0, 0,
  5.37323, _,
  0, 0,
  5.345459, _,
  0, 0,
  4.961548, _,
  0, 0,
  4.648621, _,
  0, 0,
  4.233215, _,
  0, 0,
  3.85791, _,
  0, 0,
  3.543701, _,
  0, 0,
  3.268311, _,
  0, 0,
  3.055176, _,
  0, 0,
  2.810852, _,
  0, 0,
  2.613647, _,
  0, 0,
  2.467224, _,
  0, 0,
  2.357178, _,
  0, 0,
  2.241028, _,
  0, 0,
  2.119263, _,
  0, 0,
  2.003784, _,
  0, 0,
  1.905823, _,
  0, 0,
  1.837219, _,
  0, 0,
  1.849548, _,
  0, 0,
  2.064758, _,
  0, 0,
  2.04364, _,
  0, 0,
  1.898865, _,
  0, 0,
  1.80603, _,
  0, 0,
  1.769531, _,
  0, 0,
  2.244812, _,
  0, 0,
  3.739014, _,
  0, 0,
  4.359314, _,
  0, 0,
  5.059937, _,
  0, 0,
  4.111328, _,
  0, 0,
  3.435059, _,
  0, 0,
  2.973877, _,
  0, 0,
  2.756592, _,
  0, 0,
  3.737366, _,
  0, 0,
  5.927612, _,
  0, 0,
  18.45728, _,
  0, 0,
  21.96429, _,
  0, 0,
  18.4834, _,
  0, 0,
  15.13452, _,
  0, 0,
  12.17938, _,
  0, 0,
  9.723511, _,
  0, 0,
  7.596313, _,
  0, 0,
  5.949768, _,
  0, 0,
  5.113647, _,
  0, 0,
  4.855225, _,
  0, 0,
  3.830261, _,
  0, 0,
  3.113159, _,
  0, 0,
  2.608215, _,
  0, 0,
  2.226868, _,
  0, 0,
  1.93927, _,
  0, 0,
  1.772217, _,
  0, 0,
  2.394958, _,
  0, 0,
  2.375671, _,
  0, 0,
  2.093811, _,
  0, 0,
  1.857361, _,
  0, 0,
  1.679993, _,
  0, 0,
  1.557129, _,
  0, 0,
  1.46637, _,
  0, 0,
  1.398987, _,
  0, 0,
  1.354492, _,
  0, 0,
  1.319092, _,
  0, 0,
  1.288269, _,
  0, 0,
  1.273376, _,
  0, 0,
  1.299805, _,
  0, 0,
  1.266296, _,
  0, 0,
  1.238953, _,
  0, 0,
  1.214539, _,
  0, 0,
  1.194031, _,
  0, 0,
  1.174377, _,
  0, 0,
  1.156555, _,
  0, 0,
  1.14093, _,
  0, 0,
  1.126892, _,
  0, 0,
  1.109924, _,
  0, 0,
  1.091919, _,
  0, 0,
  1.077942, _,
  0, 0,
  1.099854, _,
  0, 0,
  1.084412, _,
  0, 0,
  1.083435, _,
  0, 0,
  1.159241, _,
  0, 0,
  1.36261, _,
  0, 0,
  1.281311, _,
  0, 0,
  1.198486, _,
  0, 0,
  1.134888, _,
  0, 0,
  1.110901, _,
  0, 0,
  1.232788, _,
  0, 0,
  1.215332, _,
  0, 0,
  1.158325, _,
  0, 0,
  1.114075, _,
  0, 0,
  1.204102, _,
  0, 0,
  1.234497, _,
  0, 0,
  1.205322, _,
  0, 0,
  1.163574, _,
  0, 0,
  1.146606, _,
  0, 0,
  1.112061, _,
  0, 0,
  1.071289, _,
  0, 0,
  1.034851, _,
  0, 0,
  1.008118, _,
  0, 0,
  0.9853516, _,
  0, 0,
  0.9793701, _,
  0, 0,
  0.9710083, _,
  0, 0,
  1.136658, _,
  0, 0,
  1.408875, _,
  0, 0,
  1.376526, _,
  0, 0,
  1.300354, _,
  0, 0,
  1.817139, _,
  0, 0,
  1.893311, _,
  0, 0,
  1.780457, _,
  0, 0,
  1.652649, _,
  0, 0,
  1.546326, _,
  0, 0,
  1.456726, _,
  0, 0,
  1.374268, _,
  0, 0,
  1.305786, _,
  0, 0,
  1.251587, _,
  0, 0,
  1.201416, _,
  0, 0,
  1.158142, _,
  0, 0,
  1.13092, _,
  0, 0,
  1.24469, _,
  0, 0,
  1.309021, _,
  0, 0,
  1.266418, _,
  0, 0,
  1.223694, _,
  0, 0,
  1.180542, _,
  0, 0,
  1.139221, _,
  0, 0,
  1.101807, _,
  0, 0,
  1.070557, _,
  0, 0,
  1.045654, _,
  0, 0,
  1.040649, _,
  0, 0,
  1.064575, _,
  0, 0,
  1.045959, _,
  0, 0,
  1.071106, _,
  0, 0,
  1.362305, _,
  0, 0,
  1.448975, _,
  0, 0,
  1.43335, _,
  0, 0,
  1.424866, _,
  0, 0,
  1.545166, _,
  0, 0,
  1.527344, _,
  0, 0,
  1.463196, _,
  0, 0,
  1.429016, _,
  0, 0,
  1.428528, _,
  0, 0,
  1.400879, _,
  0, 0,
  1.392151, _,
  0, 0,
  1.662048, _,
  0, 0,
  2.14386, _,
  0, 0,
  2.224365, _,
  0, 0,
  2.143494, _,
  0, 0,
  2.083496, _,
  0, 0,
  1.998718, _,
  0, 0,
  1.912354, _,
  0, 0,
  1.833801, _,
  0, 0,
  1.75708, _,
  0, 0,
  1.686707, _,
  0, 0,
  1.639038, _,
  0, 0,
  1.578247, _,
  0, 0,
  1.53064, _,
  0, 0,
  3.261902, _,
  0, 0,
  8.547485, _,
  0, 0,
  10.51025, _,
  0, 0,
  10.26746, _,
  0, 0,
  9.740112, _,
  0, 0,
  9.254272, _,
  0, 0,
  8.725586, _,
  0, 0,
  8.156128, _,
  0, 0,
  7.517822, _,
  0, 0,
  6.955688, _,
  0, 0,
  6.5625, _,
  0, 0,
  7.245178, _,
  0, 0,
  7.048523, _,
  0, 0,
  6.536743, _,
  0, 0,
  6.167297, _,
  0, 0,
  5.848328, _,
  0, 0,
  5.658875, _,
  0, 0,
  5.88678, _,
  0, 0,
  6.60907, _,
  0, 0,
  12.25354, _,
  0, 0,
  22.29938, _,
  0, 0,
  21.42517, _,
  0, 0,
  20.58472, _,
  0, 0,
  19.72565, _,
  0, 0,
  19.19397, _,
  0, 0,
  18.70123, _,
  0, 0,
  18.09857, _,
  0, 0,
  17.53845, _,
  0, 0,
  17.08032, _,
  0, 0,
  16.60638, _,
  0, 0,
  16.03174, _,
  0, 0,
  15.58636, _,
  0, 0,
  15.91577, _,
  0, 0,
  17.9726, _,
  0, 0,
  17.75342, _,
  0, 0,
  17.11896, _,
  0, 0,
  16.5885, _,
  0, 0,
  16.42993, _,
  0, 0,
  17.10767, _,
  0, 0,
  16.38165, _,
  0, 0,
  15.82361, _,
  0, 0,
  15.40399, _,
  0, 0,
  15.16327, _,
  0, 0,
  17.31525, _,
  0, 0,
  17.17822, _,
  0, 0,
  17.82666, _,
  0, 0,
  21.54431, _,
  0, 0,
  23.86835, _,
  0, 0,
  25.3053, _,
  0, 0,
  24.23358, _,
  0, 0,
  22.604, _,
  0, 0,
  21.89081, _,
  0, 0,
  21.43756, _,
  0, 0,
  20.9115, _,
  0, 0,
  20.29425, _,
  0, 0,
  19.70282, _,
  0, 0,
  19.65503, _,
  0, 0,
  23.41473, _,
  0, 0,
  25.71649, _,
  0, 0,
  24.32574, _,
  0, 0,
  23.61914, _,
  0, 0,
  23.96582, _,
  0, 0,
  23.51898, _,
  0, 0,
  23.70404, _,
  0, 0,
  27.41412, _,
  0, 0,
  26.17462, _,
  0, 0,
  25.39343, _,
  0, 0,
  25.23944, _,
  0, 0,
  24.60791, _,
  0, 0,
  24.02783, _,
  0, 0,
  25.70483, _,
  0, 0,
  24.52222, _,
  0, 0,
  23.83484, _,
  0, 0,
  23.25635, _,
  0, 0,
  22.48804, _,
  0, 0,
  21.94775, _,
  0, 0,
  21.31226, _,
  0, 0,
  20.71484, _,
  0, 0,
  20.29578, _,
  0, 0,
  20.25354, _,
  0, 0,
  20.07751, _,
  0, 0,
  19.80621, _,
  0, 0,
  19.51331, _,
  0, 0,
  19.25244, _,
  0, 0,
  18.97815, _,
  0, 0,
  18.52991, _,
  0, 0,
  18.97833, _,
  0, 0,
  19.92194, _,
  0, 0,
  19.17902, _,
  0, 0,
  18.72394, _,
  0, 0,
  20.65369, _,
  0, 0,
  20.30286, _,
  0, 0,
  19.51697, _,
  0, 0,
  18.88147, _,
  0, 0,
  18.3891, _,
  0, 0,
  17.91058, _,
  0, 0,
  17.30426, _,
  0, 0,
  16.80072, _,
  0, 0,
  16.37537, _,
  0, 0,
  15.7793, _,
  0, 0,
  14.92328, _,
  0, 0,
  13.78894, _,
  0, 0,
  12.8537, _,
  0, 0,
  12.16064, _,
  0, 0,
  11.51111, _,
  0, 0,
  10.89117, _,
  0, 0,
  10.42767, _,
  0, 0,
  9.999695, _,
  0, 0,
  9.555786, _,
  0, 0,
  9.192505, _,
  0, 0,
  8.788391, _,
  0, 0,
  8.300964, _,
  0, 0,
  7.838867, _,
  0, 0,
  8.147278, _,
  0, 0,
  8.384277, _,
  0, 0,
  7.999878, _,
  0, 0,
  7.524231, _,
  0, 0,
  7.083496, _,
  0, 0,
  6.565918, _,
  0, 0,
  6.03656, _,
  0, 0,
  5.510803, _,
  0, 0,
  5.043091, _,
  0, 0,
  4.653381, _,
  0, 0,
  4.286377, _,
  0, 0,
  4.006775, _,
  0, 0,
  3.787231, _,
  0, 0,
  3.58905, _,
  0, 0,
  3.393494, _,
  0, 0,
  3.205017, _,
  0, 0,
  3.052002, _,
  0, 0,
  2.910828, _,
  0, 0,
  2.780029, _,
  0, 0,
  2.695679, _,
  0, 0,
  2.597107, _,
  0, 0,
  2.506836, _,
  0, 0,
  2.419983, _,
  0, 0,
  2.341675, _,
  0, 0,
  2.281799, _,
  0, 0,
  2.214478, _,
  0, 0,
  2.151855, _,
  0, 0,
  2.093262, _,
  0, 0,
  2.040405, _,
  0, 0,
  2.008057, _,
  0, 0,
  2.037659, _,
  0, 0,
  2.030457, _,
  0, 0,
  2.030945, _,
  0, 0,
  2.116333, _,
  0, 0,
  2.192505, _,
  0, 0,
  2.165466, _,
  0, 0,
  2.13446, _,
  0, 0,
  2.105713, _,
  0, 0,
  2.071594, _,
  0, 0,
  2.029053, _,
  0, 0,
  1.990173, _,
  0, 0,
  2.516479, _,
  0, 0,
  3.360168, _,
  0, 0,
  3.209473, _,
  0, 0,
  3.127197, _,
  0, 0,
  2.995667, _,
  0, 0,
  2.84259, _,
  0, 0,
  2.66272, _,
  0, 0,
  2.495483, _,
  0, 0,
  2.342285, _,
  0, 0,
  2.223267, _,
  0, 0,
  2.208374, _,
  0, 0,
  2.416931, _,
  0, 0,
  2.356018, _,
  0, 0,
  2.263611, _,
  0, 0,
  2.167847, _,
  0, 0,
  2.070984, _,
  0, 0,
  1.970276, _,
  0, 0,
  1.871765, _,
  0, 0,
  1.800232, _,
  0, 0,
  1.749451, _,
  0, 0,
  1.889038, _,
  0, 0,
  1.880615, _,
  0, 0,
  1.813965, _,
  0, 0,
  1.756042, _,
  0, 0,
  1.703308, _,
  0, 0,
  1.641663, _,
  0, 0,
  1.590027, _,
  0, 0,
  1.559326, _,
  0, 0,
  1.534485, _,
  0, 0,
  1.506226, _,
  0, 0,
  1.619019, _,
  0, 0,
  2.018433, _,
  0, 0,
  1.914429, _,
  0, 0,
  1.81488, _,
  0, 0,
  1.747009, _,
  0, 0,
  1.682251, _,
  0, 0,
  1.629761, _,
  0, 0,
  1.590149, _,
  0, 0,
  1.560608, _,
  0, 0,
  1.645386, _,
  0, 0,
  3.416687, _,
  0, 0,
  5.968262, _,
  0, 0,
  5.80658, _,
  0, 0,
  5.331421, _,
  0, 0,
  4.97406, _,
  0, 0,
  4.495972, _,
  0, 0,
  3.935913, _,
  0, 0,
  3.443054, _,
  0, 0,
  3.045044, _,
  0, 0,
  2.831421, _,
  0, 0,
  2.65564, _,
  0, 0,
  2.465637, _,
  0, 0,
  2.280945, _,
  0, 0,
  2.113953, _,
  0, 0,
  1.965698, _,
  0, 0,
  1.927185, _,
  0, 0,
  1.900513, _,
  0, 0,
  1.80188, _,
  0, 0,
  1.712036, _,
  0, 0,
  1.612061, _,
  0, 0,
  1.510071, _,
  0, 0,
  1.425598, _,
  0, 0,
  1.728088, _,
  0, 0,
  9.063354, _,
  0, 0,
  11.664, _,
  0, 0,
  9.746033, _,
  0, 0,
  8.126526, _,
  0, 0,
  6.889771, _,
  0, 0,
  5.873657, _,
  0, 0,
  5.367737, _,
  0, 0,
  5.029175, _,
  0, 0,
  4.250854, _,
  0, 0,
  4.101807, _,
  0, 0,
  5.754822, _,
  0, 0,
  5.387512, _,
  0, 0,
  4.63623, _,
  0, 0,
  7.535095, _,
  0, 0,
  11.96851, _,
  0, 0,
  10.50635, _,
  0, 0,
  9.015686, _,
  0, 0,
  7.366516, _,
  0, 0,
  6.483887, _,
  0, 0,
  6.710999, _,
  0, 0,
  6.562683, _,
  0, 0,
  6.249451, _,
  0, 0,
  6.093811, _,
  0, 0,
  4.985657, _,
  0, 0,
  4.109253, _,
  0, 0,
  3.499756, _,
  0, 0,
  3.065369, _,
  0, 0,
  2.696411, _,
  0, 0,
  2.408875, _,
  0, 0,
  2.166077, _,
  0, 0,
  1.961426, _,
  0, 0,
  1.807678, _,
  0, 0,
  1.679016, _,
  0, 0,
  1.715027, _,
  0, 0,
  1.69873, _,
  0, 0,
  2.07782, _,
  0, 0,
  3.670105, _,
  0, 0,
  4.15387, _,
  0, 0,
  3.64563, _,
  0, 0,
  3.099243, _,
  0, 0,
  2.684998, _,
  0, 0,
  2.352173, _,
  0, 0,
  2.166992, _,
  0, 0,
  1.963989, _,
  0, 0,
  1.803955, _,
  0, 0,
  1.638306, _,
  0, 0,
  1.476135, _,
  0, 0,
  1.340881, _,
  0, 0,
  1.245605, _,
  0, 0,
  1.177551, _,
  0, 0,
  1.113586, _,
  0, 0,
  1.066223, _,
  0, 0,
  1.031189, _,
  0, 0,
  0.9885254, _,
  0, 0,
  0.9510498, _,
  0, 0,
  0.9243164, _,
  0, 0,
  0.8998413, _,
  0, 0,
  0.8999023, _,
  0, 0,
  0.9855347, _,
  0, 0,
  0.9790039, _,
  0, 0,
  0.9503784, _,
  0, 0,
  0.9268799, _,
  0, 0,
  0.9046631, _,
  0, 0,
  0.8887329, _,
  0, 0,
  0.9606934, _,
  0, 0,
  0.9711914, _,
  0, 0,
  0.9414673, _,
  0, 0,
  1.234802, _,
  0, 0,
  1.854309, _,
  0, 0,
  1.829041, _,
  0, 0,
  1.692871, _,
  0, 0,
  2.502197, _,
  0, 0,
  4.354309, _,
  0, 0,
  3.684265, _,
  0, 0,
  3.135193, _,
  0, 0,
  2.692505, _,
  0, 0,
  2.340149, _,
  0, 0,
  2.053223, _,
  0, 0,
  1.942932, _,
  0, 0,
  1.794495, _,
  0, 0,
  1.643005, _,
  0, 0,
  1.523071, _,
  0, 0,
  1.423218, _,
  0, 0,
  1.32196, _,
  0, 0,
  1.233093, _,
  0, 0,
  1.160767, _,
  0, 0,
  1.09906, _,
  0, 0,
  1.047913, _,
  0, 0,
  1.013123, _,
  0, 0,
  0.9860229, _,
  0, 0,
  0.9581299, _,
  0, 0,
  0.9284058, _,
  0, 0,
  0.9005737, _,
  0, 0,
  0.8768921, _,
  0, 0,
  0.8568115, _,
  0, 0,
  0.8550415, _,
  0, 0,
  0.8479004, _,
  0, 0,
  0.8372192, _,
  0, 0,
  0.8277588, _,
  0, 0,
  0.8168945, _,
  0, 0,
  0.8058472, _,
  0, 0,
  0.7969971, _,
  0, 0,
  0.791687, _,
  0, 0,
  0.7890015, _,
  0, 0,
  0.7879028, _,
  0, 0,
  0.8861084, _,
  0, 0,
  0.9006348, _,
  0, 0,
  0.8793335, _,
  0, 0,
  0.8626099, _,
  0, 0,
  0.8496704, _,
  0, 0,
  0.8421021, _,
  0, 0,
  0.8497925, _,
  0, 0,
  0.8927612, _,
  0, 0,
  0.9348145, _,
  0, 0,
  0.928772, _,
  0, 0,
  0.9078369, _,
  0, 0,
  0.8904419, _,
  0, 0,
  0.8796387, _,
  0, 0,
  0.9521484, _,
  0, 0,
  0.9570923, _,
  0, 0,
  0.9391479, _,
  0, 0,
  0.9240112, _,
  0, 0,
  0.93573, _,
  0, 0,
  0.9256592, _,
  0, 0,
  0.9381714, _,
  0, 0,
  0.9499512, _,
  0, 0,
  0.9382935, _,
  0, 0,
  0.9261475, _,
  0, 0,
  0.9140015, _,
  0, 0,
  0.9174194, _,
  0, 0,
  0.9188232, _,
  0, 0,
  0.9254761, _,
  0, 0,
  0.9644165, _,
  0, 0,
  1.248169, _,
  0, 0,
  1.417542, _,
  0, 0,
  3.205017, _,
  0, 0,
  4.864136, _,
  0, 0,
  5.098328, _,
  0, 0,
  5.317261, _,
  0, 0,
  5.434753, _,
  0, 0,
  5.255798, _,
  0, 0,
  5.135498, _,
  0, 0,
  7.126831, _,
  0, 0,
  8.720581, _,
  0, 0,
  8.34491, _,
  0, 0,
  7.714417, _,
  0, 0,
  7.421692, _,
  0, 0,
  8.462708, _,
  0, 0,
  9.299194, _,
  0, 0,
  9.000183, _,
  0, 0,
  8.594421, _,
  0, 0,
  8.030457, _,
  0, 0,
  7.46936, _,
  0, 0,
  6.92926, _,
  0, 0,
  6.597168, _,
  0, 0,
  6.296204, _,
  0, 0,
  5.953186, _,
  0, 0,
  5.593262, _,
  0, 0,
  6.579712, _,
  0, 0,
  11.38647, _,
  0, 0,
  10.93634, _,
  0, 0,
  10.36005, _,
  0, 0,
  9.787292, _,
  0, 0,
  9.266418, _,
  0, 0,
  8.878723, _,
  0, 0,
  8.538147, _,
  0, 0,
  8.085144, _,
  0, 0,
  7.632202, _,
  0, 0,
  7.209351, _,
  0, 0,
  6.819763, _,
  0, 0,
  6.695129, _,
  0, 0,
  6.759705, _,
  0, 0,
  6.591919, _,
  0, 0,
  6.318665, _,
  0, 0,
  6.055725, _,
  0, 0,
  5.792725, _,
  0, 0,
  5.580688, _,
  0, 0,
  5.414856, _,
  0, 0,
  5.208435, _,
  0, 0,
  5.094238, _,
  0, 0,
  6.981323, _,
  0, 0,
  7.529785, _,
  0, 0,
  8.097351, _,
  0, 0,
  8.616943, _,
  0, 0,
  11.26495, _,
  0, 0,
  13.45441, _,
  0, 0,
  13.59778, _,
  0, 0,
  13.30365, _,
  0, 0,
  13.03131, _,
  0, 0,
  12.79565, _,
  0, 0,
  12.41815, _,
  0, 0,
  12.18402, _,
  0, 0,
  11.87567, _,
  0, 0,
  19.32483, _,
  0, 0,
  19.3772, _,
  0, 0,
  19.83978, _,
  0, 0,
  19.55377, _,
  0, 0,
  18.57806, _,
  0, 0,
  18.35693, _,
  0, 0,
  20.64734, _,
  0, 0,
  20.18243, _,
  0, 0,
  20.09979, _,
  0, 0,
  20.93146, _,
  0, 0,
  20.71033, _,
  0, 0,
  20.78217, _,
  0, 0,
  20.67358, _,
  0, 0,
  22.2204, _,
  0, 0,
  22.39191, _,
  0, 0,
  25.08282, _,
  0, 0,
  24.39771, _,
  0, 0,
  22.99036, _,
  0, 0,
  22.52069, _,
  0, 0,
  21.78912, _,
  0, 0,
  21.10516, _,
  0, 0,
  20.56836, _,
  0, 0,
  20.72845, _,
  0, 0,
  20.62915, _,
  0, 0,
  20.17883, _,
  0, 0,
  19.6944, _,
  0, 0,
  19.46021, _,
  0, 0,
  18.91309, _,
  0, 0,
  18.17535, _,
  0, 0,
  17.65314, _,
  0, 0,
  17.12738, _,
  0, 0,
  18.164, _,
  0, 0,
  21.37354, _,
  0, 0,
  23.03265, _,
  0, 0,
  27.13983, _,
  0, 0,
  24.78595, _,
  0, 0,
  23.67725, _,
  0, 0,
  23.02393, _,
  0, 0,
  22.4223, _,
  0, 0,
  23.20312, _,
  0, 0,
  23.44904, _,
  0, 0,
  24.70935, _,
  0, 0,
  23.62524, _,
  0, 0,
  24.33136, _,
  0, 0,
  24.01123, _,
  0, 0,
  23.24097, _,
  0, 0,
  22.58478, _,
  0, 0,
  21.91553, _,
  0, 0,
  21.45959, _,
  0, 0,
  21.02466, _,
  0, 0,
  20.34705, _,
  0, 0,
  20.659, _,
  0, 0,
  21.67633, _,
  0, 0,
  20.89221, _,
  0, 0,
  20.16766, _,
  0, 0,
  19.42688, _,
  0, 0,
  18.76135, _,
  0, 0,
  18.08014, _,
  0, 0,
  17.27209, _,
  0, 0,
  16.49365, _,
  0, 0,
  15.74097, _,
  0, 0,
  15.82776, _,
  0, 0,
  16.25684, _,
  0, 0,
  15.68463, _,
  0, 0,
  14.99719, _,
  0, 0,
  14.28119, _,
  0, 0,
  13.5282, _,
  0, 0,
  12.89136, _,
  0, 0,
  12.27692, _,
  0, 0,
  11.99139, _,
  0, 0,
  11.97101, _,
  0, 0,
  11.51245, _,
  0, 0,
  10.78485, _,
  0, 0,
  10.01263, _,
  0, 0,
  9.238464, _,
  0, 0,
  8.449219, _,
  0, 0,
  8.34375, _,
  0, 0,
  8.329712, _,
  0, 0,
  7.894165, _,
  0, 0,
  7.319946, _,
  0, 0,
  6.829895, _,
  0, 0,
  6.340942, _,
  0, 0,
  6.033203, _,
  0, 0,
  5.69574, _,
  0, 0,
  8.908203, _,
  0, 0,
  12.59448, _,
  0, 0,
  14.17151, _,
  0, 0,
  14.23145, _,
  0, 0,
  13.64856, _,
  0, 0,
  12.83154, _,
  0, 0,
  11.76538, _,
  0, 0,
  10.66833, _,
  0, 0,
  9.602234, _,
  0, 0,
  8.614319, _,
  0, 0,
  7.690735, _,
  0, 0,
  6.835815, _,
  0, 0,
  6.091187, _,
  0, 0,
  5.575317, _,
  0, 0,
  5.361206, _,
  0, 0,
  5.103821, _,
  0, 0,
  5.989502, _,
  0, 0,
  6.046631, _,
  0, 0,
  9.329346, _,
  0, 0,
  11.51819, _,
  0, 0,
  13.58875, _,
  0, 0,
  12.91412, _,
  0, 0,
  13.22345, _,
  0, 0,
  13.25818, _,
  0, 0,
  13.89093, _,
  0, 0,
  13.18951, _,
  0, 0,
  13.65839, _,
  0, 0,
  14.29211, _,
  0, 0,
  16.55835, _,
  0, 0,
  15.22058, _,
  0, 0,
  13.50104, _,
  0, 0,
  11.77216, _,
  0, 0,
  11.28235, _,
  0, 0,
  10.38153, _,
  0, 0,
  9.092407, _,
  0, 0,
  7.857422, _,
  0, 0,
  6.72229, _,
  0, 0,
  5.733704, _,
  0, 0,
  4.88147, _,
  0, 0,
  4.197327, _,
  0, 0,
  3.660889, _,
  0, 0,
  3.246704, _,
  0, 0,
  2.914734, _,
  0, 0,
  2.651978, _,
  0, 0,
  2.398132, _,
  0, 0,
  2.196411, _,
  0, 0,
  3.883728, _,
  0, 0,
  5.147766, _,
  0, 0,
  4.812561, _,
  0, 0,
  4.66095, _,
  0, 0,
  4.288208, _,
  0, 0,
  3.81311, _,
  0, 0,
  3.382812, _,
  0, 0,
  3.591309, _,
  0, 0,
  14.24481, _,
  0, 0,
  28.4516, _,
  0, 0,
  29.73926, _,
  0, 0,
  27.16339, _,
  0, 0,
  24.81775, _,
  0, 0,
  22.49756, _,
  0, 0,
  19.80322, _,
  0, 0,
  17.85333, _,
  0, 0,
  16.01282, _,
  0, 0,
  14.07953, _,
  0, 0,
  11.95526, _,
  0, 0,
  10.05524, _,
  0, 0,
  8.431213, _,
  0, 0,
  7.0495, _,
  0, 0,
  5.879089, _,
  0, 0,
  4.922668, _,
  0, 0,
  4.164673, _,
  0, 0,
  3.659302, _,
  0, 0,
  3.350525, _,
  0, 0,
  3.112793, _,
  0, 0,
  3.014587, _,
  0, 0,
  2.858276, _,
  0, 0,
  2.787292, _,
  0, 0,
  2.633362, _,
  0, 0,
  2.587952, _,
  0, 0,
  2.696411, _,
  0, 0,
  2.523621, _,
  0, 0,
  2.359558, _,
  0, 0,
  2.721436, _,
  0, 0,
  2.962891, _,
  0, 0,
  3.039917, _,
  0, 0,
  2.90509, _,
  0, 0,
  2.641357, _,
  0, 0,
  2.369812, _,
  0, 0,
  2.231995, _,
  0, 0,
  2.232544, _,
  0, 0,
  2.264404, _,
  0, 0,
  2.132446, _,
  0, 0,
  2.129822, _,
  0, 0,
  4.845886, _,
  0, 0,
  4.773132, _,
  0, 0,
  4.169128, _,
  0, 0,
  3.639465, _,
  0, 0,
  3.203247, _,
  0, 0,
  2.885071, _,
  0, 0,
  2.64679, _,
  0, 0,
  2.721619, _,
  0, 0,
  2.873779, _,
  0, 0,
  2.610657, _,
  0, 0,
  2.37738, _,
  0, 0,
  2.159241, _,
  0, 0,
  2.188965, _,
  0, 0,
  5.615662, _,
  0, 0,
  8.555908, _,
  0, 0,
  7.275757, _,
  0, 0,
  6.176208, _,
  0, 0,
  7.214966, _,
  0, 0,
  8.80127, _,
  0, 0,
  7.823853, _,
  0, 0,
  11.15869, _,
  0, 0,
  10.99548, _,
  0, 0,
  8.899597, _,
  0, 0,
  7.152161, _,
  0, 0,
  5.828369, _,
  0, 0,
  4.790222, _,
  0, 0,
  4.036804, _,
  0, 0,
  3.463562, _,
  0, 0,
  3.002319, _,
  0, 0,
  2.60553, _,
  0, 0,
  2.273743, _,
  0, 0,
  2.04657, _,
  0, 0,
  1.882751, _,
  0, 0,
  1.738159, _,
  0, 0,
  1.606873, _,
  0, 0,
  1.493408, _,
  0, 0,
  1.394409, _,
  0, 0,
  1.324951, _,
  0, 0,
  1.269836, _,
  0, 0,
  1.227356, _,
  0, 0,
  1.242859, _,
  0, 0,
  1.210449, _,
  0, 0,
  1.169739, _,
  0, 0,
  1.138245, _,
  0, 0,
  1.197937, _,
  0, 0,
  1.208069, _,
  0, 0,
  1.177124, _,
  0, 0,
  1.147644, _,
  0, 0,
  1.122803, _,
  0, 0,
  1.100098, _,
  0, 0,
  1.08075, _,
  0, 0,
  1.059509, _,
  0, 0,
  1.040222, _,
  0, 0,
  1.027039, _,
  0, 0,
  1.015686, _,
  0, 0,
  1.004395, _,
  0, 0,
  0.9917603, _,
  0, 0,
  0.982666, _,
  0, 0,
  0.9793091, _,
  0, 0,
  0.9755859, _,
  0, 0,
  0.9691162, _,
  0, 0,
  0.9606323, _,
  0, 0,
  0.9524536, _,
  0, 0,
  0.9455566, _,
  0, 0,
  0.9377441, _,
  0, 0,
  0.9312744, _,
  0, 0,
  0.9255371, _,
  0, 0,
  0.9194946, _,
  0, 0,
  0.9107666, _,
  0, 0,
  0.9002075, _,
  0, 0,
  0.8937988, _,
  0, 0,
  0.8912354, _,
  0, 0,
  0.8889771, _,
  0, 0,
  0.8849487, _,
  0, 0,
  0.8796997, _,
  0, 0,
  0.8753052, _,
  0, 0,
  0.8770752, _,
  0, 0,
  0.8894043, _,
  0, 0,
  0.9058838, _,
  0, 0,
  1.010071, _,
  0, 0,
  1.119141, _,
  0, 0,
  1.079285, _,
  0, 0,
  1.031921, _,
  0, 0,
  0.9920044, _,
  0, 0,
  1.035461, _,
  0, 0,
  1.25238, _,
  0, 0,
  1.653076, _,
  0, 0,
  1.968445, _,
  0, 0,
  2.16803, _,
  0, 0,
  2.657593, _,
  0, 0,
  2.772827, _,
  0, 0,
  2.614807, _,
  0, 0,
  5.355164, _,
  0, 0,
  7.196228, _,
  0, 0,
  7.105896, _,
  0, 0,
  7.047485, _,
  0, 0,
  10.17456, _,
  0, 0,
  11.27563, _,
  0, 0,
  9.789124, _,
  0, 0,
  8.493408, _,
  0, 0,
  7.57605, _,
  0, 0,
  7.089417, _,
  0, 0,
  7.19696, _,
  0, 0,
  9.223877, _,
  0, 0,
  10.20508, _,
  0, 0,
  9.023804, _,
  0, 0,
  8.02887, _,
  0, 0,
  7.231323, _,
  0, 0,
  12.76172, _,
  0, 0,
  14.99243, _,
  0, 0,
  22.44196, _,
  0, 0,
  21.19635, _,
  0, 0,
  18.84607, _,
  0, 0,
  16.88745, _,
  0, 0,
  14.98877, _,
  0, 0,
  13.38916, _,
  0, 0,
  11.94543, _,
  0, 0,
  10.79614, _,
  0, 0,
  9.908752, _,
  0, 0,
  10.4754, _,
  0, 0,
  12.68097, _,
  0, 0,
  12.76556, _,
  0, 0,
  11.76904, _,
  0, 0,
  10.75037, _,
  0, 0,
  10.5993, _,
  0, 0,
  11.60535, _,
  0, 0,
  16.383, _,
  0, 0,
  20.03125, _,
  0, 0,
  20.43384, _,
  0, 0,
  19.32428, _,
  0, 0,
  18.5528, _,
  0, 0,
  17.56146, _,
  0, 0,
  16.64551, _,
  0, 0,
  16.45026, _,
  0, 0,
  15.86481, _,
  0, 0,
  15.06927, _,
  0, 0,
  14.35284, _,
  0, 0,
  13.23663, _,
  0, 0,
  12.1662, _,
  0, 0,
  11.99402, _,
  0, 0,
  13.66095, _,
  0, 0,
  18.6015, _,
  0, 0,
  17.83453, _,
  0, 0,
  16.93256, _,
  0, 0,
  15.91284, _,
  0, 0,
  14.94806, _,
  0, 0,
  14.04572, _,
  0, 0,
  12.97314, _,
  0, 0,
  11.75281, _,
  0, 0,
  10.8244, _,
  0, 0,
  10.23596, _,
  0, 0,
  9.731323, _,
  0, 0,
  9.36377, _,
  0, 0,
  9.045471, _,
  0, 0,
  8.619263, _,
  0, 0,
  8.277344, _,
  0, 0,
  7.946655, _,
  0, 0,
  7.586121, _,
  0, 0,
  7.381348, _,
  0, 0,
  7.143982, _,
  0, 0,
  6.848145, _,
  0, 0,
  6.795654, _,
  0, 0,
  6.639648, _,
  0, 0,
  6.556824, _,
  0, 0,
  6.424561, _,
  0, 0,
  7.025452, _,
  0, 0,
  7.002319, _,
  0, 0,
  6.663086, _,
  0, 0,
  10.43341, _,
  0, 0,
  17.10455, _,
  0, 0,
  17.69812, _,
  0, 0,
  17.27405, _,
  0, 0,
  17.9386, _,
  0, 0,
  18.42102, _,
  0, 0,
  18.06506, _,
  0, 0,
  17.63025, _,
  0, 0,
  17.08972, _,
  0, 0,
  16.65845, _,
  0, 0,
  16.53125, _,
  0, 0,
  15.89294, _,
  0, 0,
  17.71252, _,
  0, 0,
  19.87775, _,
  0, 0,
  19.31818, _,
  0, 0,
  18.57965, _,
  0, 0,
  18.0022, _,
  0, 0,
  17.51611, _,
  0, 0,
  17.11847, _,
  0, 0,
  17.77826, _,
  0, 0,
  17.68176, _,
  0, 0,
  17.09247, _,
  0, 0,
  16.45532, _,
  0, 0,
  15.84906, _,
  0, 0,
  16.22491, _,
  0, 0,
  16.45349, _,
  0, 0,
  16.01202, _,
  0, 0,
  15.4884, _,
  0, 0,
  14.89636, _,
  0, 0,
  15.0473, _,
  0, 0,
  14.59119, _,
  0, 0,
  13.98981, _,
  0, 0,
  13.46686, _,
  0, 0,
  13.03619, _,
  0, 0,
  12.66388, _,
  0, 0,
  12.31061, _,
  0, 0,
  11.98895, _,
  0, 0,
  11.75494, _,
  0, 0,
  11.43677, _,
  0, 0,
  11.12854, _,
  0, 0,
  14.1795, _,
  0, 0,
  15.13403, _,
  0, 0,
  14.70728, _,
  0, 0,
  14.31781, _,
  0, 0,
  14.19421, _,
  0, 0,
  14.18927, _,
  0, 0,
  14.28888, _,
  0, 0,
  14.23572, _,
  0, 0,
  14.08655, _,
  0, 0,
  14.07776, _,
  0, 0,
  14.09155, _,
  0, 0,
  14.69165, _,
  0, 0,
  15.9975, _,
  0, 0,
  15.74457, _,
  0, 0,
  15.28387, _,
  0, 0,
  14.7489, _,
  0, 0,
  14.1817, _,
  0, 0,
  13.61005, _,
  0, 0,
  13.02277, _,
  0, 0,
  12.44067, _,
  0, 0,
  11.95386, _,
  0, 0,
  11.61072, _,
  0, 0,
  13.80219, _,
  0, 0,
  13.53265, _,
  0, 0,
  12.97784, _,
  0, 0,
  12.21613, _,
  0, 0,
  11.638, _,
  0, 0,
  12.1651, _,
  0, 0,
  12.65308, _,
  0, 0,
  12.5412, _,
  0, 0,
  12.75867, _,
  0, 0,
  12.42432, _,
  0, 0,
  11.74994, _,
  0, 0,
  11.52832, _,
  0, 0,
  11.77216, _,
  0, 0,
  11.08386, _,
  0, 0,
  10.41705, _,
  0, 0,
  11.35028, _,
  0, 0,
  13.42255, _,
  0, 0,
  12.68781, _,
  0, 0,
  11.90619, _,
  0, 0,
  11.15582, _,
  0, 0,
  10.40021, _,
  0, 0,
  9.708923, _,
  0, 0,
  10.50537, _,
  0, 0,
  11.01434, _,
  0, 0,
  10.37616, _,
  0, 0,
  9.803955, _,
  0, 0,
  9.500427, _,
  0, 0,
  10.89374, _,
  0, 0,
  10.80725, _,
  0, 0,
  10.08746, _,
  0, 0,
  9.447815, _,
  0, 0,
  8.772888, _,
  0, 0,
  8.130737, _,
  0, 0,
  7.612915, _,
  0, 0,
  8.948792, _,
  0, 0,
  8.524353, _,
  0, 0,
  8.594177, _,
  0, 0,
  10.00604, _,
  0, 0,
  10.37433, _,
  0, 0,
  10.72021, _,
  0, 0,
  15.82672, _,
  0, 0,
  15.14099, _,
  0, 0,
  13.66589, _,
  0, 0,
  12.00854, _,
  0, 0,
  10.87634, _,
  0, 0,
  20.00183, _,
  0, 0,
  20.02576, _,
  0, 0,
  17.72015, _,
  0, 0,
  16.01233, _,
  0, 0,
  15.11829, _,
  0, 0,
  13.79773, _,
  0, 0,
  14.13684, _,
  0, 0,
  16.19806, _,
  0, 0,
  19.87567, _,
  0, 0,
  22.62085, _,
  0, 0,
  28.10944, _,
  0, 0,
  30.7207, _,
  0, 0,
  28.19409, _,
  0, 0,
  26.02057, _,
  0, 0,
  25.75592, _,
  0, 0,
  25.47479, _,
  0, 0,
  24.02399, _,
  0, 0,
  22.20105, _,
  0, 0,
  20.47986, _,
  0, 0,
  21.28546, _,
  0, 0,
  21.74597, _,
  0, 0,
  22.6001, _,
  0, 0,
  22.224, _,
  0, 0,
  22.98096, _,
  0, 0,
  22.75183, _,
  0, 0,
  20.81427, _,
  0, 0,
  19.19952, _,
  0, 0,
  17.21246, _,
  0, 0,
  15.50482, _,
  0, 0,
  13.93787, _,
  0, 0,
  12.1947, _,
  0, 0,
  10.87769, _,
  0, 0,
  11.30664, _,
  0, 0,
  11.29651, _,
  0, 0,
  9.979553, _,
  0, 0,
  9.085815, _,
  0, 0,
  9.847656, _,
  0, 0,
  10.07977, _,
  0, 0,
  9.628418, _,
  0, 0,
  9.112549, _,
  0, 0,
  8.58075, _,
  0, 0,
  7.938293, _,
  0, 0,
  7.161987, _,
  0, 0,
  6.359802, _,
  0, 0,
  5.689026, _,
  0, 0,
  5.100647, _,
  0, 0,
  4.47998, _,
  0, 0,
  3.870789, _,
  0, 0,
  3.433533, _,
  0, 0,
  3.345337, _,
  0, 0,
  3.163879, _,
  0, 0,
  2.961243, _,
  0, 0,
  2.779053, _,
  0, 0,
  2.6073, _,
  0, 0,
  2.454773, _,
  0, 0,
  2.307434, _,
  0, 0,
  2.202576, _,
  0, 0,
  2.164673, _,
  0, 0,
  5.197632, _,
  0, 0,
  5.750427, _,
  0, 0,
  6.61438, _,
  0, 0,
  7.148499, _,
  0, 0,
  6.529358, _,
  0, 0,
  6.386108, _,
  0, 0,
  5.616638, _,
  0, 0,
  4.850403, _,
  0, 0,
  4.174927, _,
  0, 0,
  3.666748, _,
  0, 0,
  4.31488, _,
  0, 0,
  4.865906, _,
  0, 0,
  4.696899, _,
  0, 0,
  4.175232, _,
  0, 0,
  3.738953, _,
  0, 0,
  3.360291, _,
  0, 0,
  3.017517, _,
  0, 0,
  2.946838, _,
  0, 0,
  2.819641, _,
  0, 0,
  3.314087, _,
  0, 0,
  3.515503, _,
  0, 0,
  3.880188, _,
  0, 0,
  3.688171, _,
  0, 0,
  3.211609, _,
  0, 0,
  2.802002, _,
  0, 0,
  2.482727, _,
  0, 0,
  2.236816, _,
  0, 0,
  2.075256, _,
  0, 0,
  1.943726, _,
  0, 0,
  1.853271, _,
  0, 0,
  1.807739, _,
  0, 0,
  1.725281, _,
  0, 0,
  1.647949, _,
  0, 0,
  1.589478, _,
  0, 0,
  1.542603, _,
  0, 0,
  1.490051, _,
  0, 0,
  1.438904, _,
  0, 0,
  1.415344, _,
  0, 0,
  1.481445, _,
  0, 0,
  1.41095, _,
  0, 0,
  1.361877, _,
  0, 0,
  1.330566, _,
  0, 0,
  1.35675, _,
  0, 0,
  1.346252, _,
  0, 0,
  1.349548, _,
  0, 0,
  1.375854, _,
  0, 0,
  1.329163, _,
  0, 0,
  1.281982, _,
  0, 0,
  1.319214, _,
  0, 0,
  1.317078, _,
  0, 0,
  1.268982, _,
  0, 0,
  1.21582, _,
  0, 0,
  1.172302, _,
  0, 0,
  1.1427, _,
  0, 0,
  1.126831, _,
  0, 0,
  1.122131, _,
  0, 0,
  1.1203, _,
  0, 0,
  1.120911, _,
  0, 0,
  1.108948, _,
  0, 0,
  1.110352, _,
  0, 0,
  1.09967, _,
  0, 0,
  1.085266, _,
  0, 0,
  1.071533, _,
  0, 0,
  1.056213, _,
  0, 0,
  1.046326, _,
  0, 0,
  1.037964, _,
  0, 0,
  1.02533, _,
  0, 0,
  1.009033, _,
  0, 0,
  0.9969482, _,
  0, 0,
  0.9862061, _,
  0, 0,
  0.9742432, _,
  0, 0,
  0.9641113, _,
  0, 0,
  0.9549561, _,
  0, 0,
  0.9481812, _,
  0, 0,
  0.9508667, _,
  0, 0,
  1.010315, _,
  0, 0,
  1.108887, _,
  0, 0,
  1.14563, _,
  0, 0,
  1.087219, _,
  0, 0,
  1.038269, _,
  0, 0,
  0.9992065, _,
  0, 0,
  0.9769287, _,
  0, 0,
  0.9656372, _,
  0, 0,
  0.9589233, _,
  0, 0,
  0.9506836, _,
  0, 0,
  0.9399414, _,
  0, 0,
  0.9272461, _,
  0, 0,
  0.9135742, _,
  0, 0,
  0.9411621, _,
  0, 0,
  0.9568481, _,
  0, 0,
  0.9330444, _,
  0, 0,
  0.9962158, _,
  0, 0,
  1.343079, _,
  0, 0,
  1.325684, _,
  0, 0,
  1.266785, _,
  0, 0,
  1.192444, _,
  0, 0,
  1.126465, _,
  0, 0,
  1.076111, _,
  0, 0,
  1.030396, _,
  0, 0,
  0.9852905, _,
  0, 0,
  1.033997, _,
  0, 0,
  1.080322, _,
  0, 0,
  1.043274, _,
  0, 0,
  1.010071, _,
  0, 0,
  0.9806519, _,
  0, 0,
  0.9933472, _,
  0, 0,
  1.132874, _,
  0, 0,
  1.125916, _,
  0, 0,
  1.406616, _,
  0, 0,
  1.457947, _,
  0, 0,
  1.583862, _,
  0, 0,
  1.94812, _,
  0, 0,
  2.096497, _,
  0, 0,
  1.977112, _,
  0, 0,
  1.815369, _,
  0, 0,
  1.68573, _,
  0, 0,
  1.582031, _,
  0, 0,
  1.512573, _,
  0, 0,
  1.512085, _,
  0, 0,
  1.676697, _,
  0, 0,
  1.952087, _,
  0, 0,
  1.893677, _,
  0, 0,
  1.799011, _,
  0, 0,
  3.789795, _,
  0, 0,
  6.170227, _,
  0, 0,
  5.309265, _,
  0, 0,
  4.72876, _,
  0, 0,
  4.279297, _,
  0, 0,
  3.836731, _,
  0, 0,
  3.479248, _,
  0, 0,
  3.197021, _,
  0, 0,
  2.954224, _,
  0, 0,
  2.821106, _,
  0, 0,
  3.087036, _,
  0, 0,
  3.269897, _,
  0, 0,
  3.439148, _,
  0, 0,
  3.340698, _,
  0, 0,
  3.962952, _,
  0, 0,
  6.64209, _,
  0, 0,
  6.843201, _,
  0, 0,
  6.077271, _,
  0, 0,
  5.627197, _,
  0, 0,
  5.92157, _,
  0, 0,
  5.898804, _,
  0, 0,
  5.791931, _,
  0, 0,
  8.365723, _,
  0, 0,
  17.23694, _,
  0, 0,
  17.25995, _,
  0, 0,
  16.11182, _,
  0, 0,
  17.91302, _,
  0, 0,
  17.7348, _,
  0, 0,
  16.66272, _,
  0, 0,
  15.65564, _,
  0, 0,
  14.43616, _,
  0, 0,
  13.30402, _,
  0, 0,
  12.60437, _,
  0, 0,
  12.20825, _,
  0, 0,
  11.8241, _,
  0, 0,
  11.15063, _,
  0, 0,
  10.21674, _,
  0, 0,
  9.222412, _,
  0, 0,
  8.098633, _,
  0, 0,
  7.125183, _,
  0, 0,
  6.703186, _,
  0, 0,
  8.922424, _,
  0, 0,
  12.47339, _,
  0, 0,
  13.49213, _,
  0, 0,
  12.46936, _,
  0, 0,
  11.4223, _,
  0, 0,
  10.5083, _,
  0, 0,
  10.24176, _,
  0, 0,
  11.30682, _,
  0, 0,
  10.66589, _,
  0, 0,
  9.949768, _,
  0, 0,
  10.48834, _,
  0, 0,
  12.36407, _,
  0, 0,
  11.71857, _,
  0, 0,
  11.07587, _,
  0, 0,
  10.52325, _,
  0, 0,
  9.974121, _,
  0, 0,
  9.372131, _,
  0, 0,
  8.815369, _,
  0, 0,
  8.338013, _,
  0, 0,
  8.561951, _,
  0, 0,
  8.868652, _,
  0, 0,
  8.490479, _,
  0, 0,
  8.968018, _,
  0, 0,
  9.28302, _,
  0, 0,
  8.873779, _,
  0, 0,
  8.419678, _,
  0, 0,
  7.947754, _,
  0, 0,
  7.464294, _,
  0, 0,
  7.288391, _,
  0, 0,
  8.479492, _,
  0, 0,
  8.251709, _,
  0, 0,
  8.437317, _,
  0, 0,
  8.455322, _,
  0, 0,
  8.969482, _,
  0, 0,
  9.545776, _,
  0, 0,
  14.62323, _,
  0, 0,
  14.47473, _,
  0, 0,
  13.995, _,
  0, 0,
  13.54498, _,
  0, 0,
  13.07849, _,
  0, 0,
  12.64606, _,
  0, 0,
  12.3222, _,
  0, 0,
  11.98627, _,
  0, 0,
  11.61627, _,
  0, 0,
  11.29584, _,
  0, 0,
  11.05066, _,
  0, 0,
  10.96912, _,
  0, 0,
  11.05035, _,
  0, 0,
  10.98523, _,
  0, 0,
  10.86658, _,
  0, 0,
  10.98254, _,
  0, 0,
  11.29156, _,
  0, 0,
  11.07605, _,
  0, 0,
  10.94641, _,
  0, 0,
  11.43225, _,
  0, 0,
  11.25677, _,
  0, 0,
  15.3855, _,
  0, 0,
  19.07056, _,
  0, 0,
  19.15088, _,
  0, 0,
  19.45514, _,
  0, 0,
  18.39447, _,
  0, 0,
  17.68585, _,
  0, 0,
  17.16003, _,
  0, 0,
  16.63953, _,
  0, 0,
  16.05762, _,
  0, 0,
  15.45813, _,
  0, 0,
  14.92938, _,
  0, 0,
  14.43085, _,
  0, 0,
  14.05554, _,
  0, 0,
  13.65283, _,
  0, 0,
  13.21783, _,
  0, 0,
  12.76447, _,
  0, 0,
  12.25183, _,
  0, 0,
  11.81128, _,
  0, 0,
  11.41077, _,
  0, 0,
  12.23956, _,
  0, 0,
  11.96069, _,
  0, 0,
  12.513, _,
  0, 0,
  12.35065, _,
  0, 0,
  12.07129, _,
  0, 0,
  12.14154, _,
  0, 0,
  13.4552, _,
  0, 0,
  13.67749, _,
  0, 0,
  13.2002, _,
  0, 0,
  12.67609, _,
  0, 0,
  12.22516, _,
  0, 0,
  11.72839, _,
  0, 0,
  11.16064, _,
  0, 0,
  10.95258, _,
  0, 0,
  11.19641, _,
  0, 0,
  11.53351, _,
  0, 0,
  11.01617, _,
  0, 0,
  10.40521, _,
  0, 0,
  9.772461, _,
  0, 0,
  9.215332, _,
  0, 0,
  9.137756, _,
  0, 0,
  8.672974, _,
  0, 0,
  8.10437, _,
  0, 0,
  7.652405, _,
  0, 0,
  7.254822, _,
  0, 0,
  6.828613, _,
  0, 0,
  6.509583, _,
  0, 0,
  6.379211, _,
  0, 0,
  6.162659, _,
  0, 0,
  5.87738, _,
  0, 0,
  5.595886, _,
  0, 0,
  5.328247, _,
  0, 0,
  5.05896, _,
  0, 0,
  4.8302, _,
  0, 0,
  4.597778, _,
  0, 0,
  4.370178, _,
  0, 0,
  4.151794, _,
  0, 0,
  4.008179, _,
  0, 0,
  3.847351, _,
  0, 0,
  3.663086, _,
  0, 0,
  3.491821, _,
  0, 0,
  3.635864, _,
  0, 0,
  3.592346, _,
  0, 0,
  3.479919, _,
  0, 0,
  3.332214, _,
  0, 0,
  3.169189, _,
  0, 0,
  3.014587, _,
  0, 0,
  2.931946, _,
  0, 0,
  3.047668, _,
  0, 0,
  3.022339, _,
  0, 0,
  2.930481, _,
  0, 0,
  2.819885, _,
  0, 0,
  2.849365, _,
  0, 0,
  3.383301, _,
  0, 0,
  6.96936, _,
  0, 0,
  7.535278, _,
  0, 0,
  6.915283, _,
  0, 0,
  6.398132, _,
  0, 0,
  5.928772, _,
  0, 0,
  6.090576, _,
  0, 0,
  5.78833, _,
  0, 0,
  5.356384, _,
  0, 0,
  4.889343, _,
  0, 0,
  4.477478, _,
  0, 0,
  4.189087, _,
  0, 0,
  3.899841, _,
  0, 0,
  9.43573, _,
  0, 0,
  11.42285, _,
  0, 0,
  11.73065, _,
  0, 0,
  11.96918, _,
  0, 0,
  10.90808, _,
  0, 0,
  9.847473, _,
  0, 0,
  9.077393, _,
  0, 0,
  8.814575, _,
  0, 0,
  8.274109, _,
  0, 0,
  7.682129, _,
  0, 0,
  7.05896, _,
  0, 0,
  7.150757, _,
  0, 0,
  7.278931, _,
  0, 0,
  6.871887, _,
  0, 0,
  7.117004, _,
  0, 0,
  6.911072, _,
  0, 0,
  12.07239, _,
  0, 0,
  16.52325, _,
  0, 0,
  14.69025, _,
  0, 0,
  13.13513, _,
  0, 0,
  11.72913, _,
  0, 0,
  10.32318, _,
  0, 0,
  9.219055, _,
  0, 0,
  8.006714, _,
  0, 0,
  7.339905, _,
  0, 0,
  12.29681, _,
  0, 0,
  12.30371, _,
  0, 0,
  10.62048, _,
  0, 0,
  9.358337, _,
  0, 0,
  8.384277, _,
  0, 0,
  7.392944, _,
  0, 0,
  6.424744, _,
  0, 0,
  5.586914, _,
  0, 0,
  4.937988, _,
  0, 0,
  4.396973, _,
  0, 0,
  3.950195, _,
  0, 0,
  3.60614, _,
  0, 0,
  3.244995, _,
  0, 0,
  2.933411, _,
  0, 0,
  2.714783, _,
  0, 0,
  2.559814, _,
  0, 0,
  2.415222, _,
  0, 0,
  2.27832, _,
  0, 0,
  2.124146, _,
  0, 0,
  2.389404, _,
  0, 0,
  10.29712, _,
  0, 0,
  14.86237, _,
  0, 0,
  15.90118, _,
  0, 0,
  15.8952, _,
  0, 0,
  14.91919, _,
  0, 0,
  15.49695, _,
  0, 0,
  16.0072, _,
  0, 0,
  14.05017, _,
  0, 0,
  11.75531, _,
  0, 0,
  9.705872, _,
  0, 0,
  7.970947, _,
  0, 0,
  9.755188, _,
  0, 0,
  9.418884, _,
  0, 0,
  7.743164, _,
  0, 0,
  6.77478, _,
  0, 0,
  8.25293, _,
  0, 0,
  7.152039, _,
  0, 0,
  6.131531, _,
  0, 0,
  5.167786, _,
  0, 0,
  4.314697, _,
  0, 0,
  3.938477, _,
  0, 0,
  3.936462, _,
  0, 0,
  3.419067, _,
  0, 0,
  3.357666, _,
  0, 0,
  3.210876, _,
  0, 0,
  2.793213, _,
  0, 0,
  2.450745, _,
  0, 0,
  2.176086, _,
  0, 0,
  2.017761, _,
  0, 0,
  1.817261, _,
  0, 0,
  1.652832, _,
  0, 0,
  1.514343, _,
  0, 0,
  1.487366, _,
  0, 0,
  2.352844, _,
  0, 0,
  3.461121, _,
  0, 0,
  3.201355, _,
  0, 0,
  3.477051, _,
  0, 0,
  4.218201, _,
  0, 0,
  5.624146, _,
  0, 0,
  4.742126, _,
  0, 0,
  4.864319, _,
  0, 0,
  4.019104, _,
  0, 0,
  3.323425, _,
  0, 0,
  3.156982, _,
  0, 0,
  2.940308, _,
  0, 0,
  2.558411, _,
  0, 0,
  2.360901, _,
  0, 0,
  2.093872, _,
  0, 0,
  1.881897, _,
  0, 0,
  1.687439, _,
  0, 0,
  1.533386, _,
  0, 0,
  1.417847, _,
  0, 0,
  1.312744, _,
  0, 0,
  1.212097, _,
  0, 0,
  1.136292, _,
  0, 0,
  1.082031, _,
  0, 0,
  1.035583, _,
  0, 0,
  0.9942627, _,
  0, 0,
  0.9578247, _,
  0, 0,
  0.928772, _,
  0, 0,
  0.9056396, _,
  0, 0,
  0.8838501, _,
  0, 0,
  0.866333, _,
  0, 0,
  0.8646851, _,
  0, 0,
  0.9150391, _,
  0, 0,
  0.9312134, _,
  0, 0,
  0.9030151, _,
  0, 0,
  0.8745728, _,
  0, 0,
  0.8521118, _,
  0, 0,
  0.8356934, _,
  0, 0,
  0.8233643, _,
  0, 0,
  0.8145752, _,
  0, 0,
  0.8088989, _,
  0, 0,
  0.8010864, _,
  0, 0,
  0.7923584, _,
  0, 0,
  0.7861938, _,
  0, 0,
  0.7813721, _,
  0, 0,
  0.7800903, _,
  0, 0,
  0.7791748, _,
  0, 0,
  0.7774658, _,
  0, 0,
  0.7745972, _,
  0, 0,
  0.7711792, _,
  0, 0,
  0.7722168, _,
  0, 0,
  0.8179321, _,
  0, 0,
  0.8182373, _,
  0, 0,
  0.80896, _,
  0, 0,
  0.7977295, _,
  0, 0,
  0.7866821, _,
  0, 0,
  0.7919312, _,
  0, 0,
  1.067261, _,
  0, 0,
  1.643372, _,
  0, 0,
  1.813232, _,
  0, 0,
  1.658569, _,
  0, 0,
  1.508423, _,
  0, 0,
  1.375977, _,
  0, 0,
  1.259338, _,
  0, 0,
  1.162659, _,
  0, 0,
  1.084045, _,
  0, 0,
  1.018372, _,
  0, 0,
  0.9640503, _,
  0, 0,
  0.9177856, _,
  0, 0,
  0.8795166, _,
  0, 0,
  0.8505859, _,
  0, 0,
  0.8253784, _,
  0, 0,
  0.8059082, _,
  0, 0,
  0.793457, _,
  0, 0,
  0.7839355, _,
  0, 0,
  0.7733765, _,
  0, 0,
  0.7658081, _,
  0, 0,
  0.7612915, _,
  0, 0,
  0.7591553, _,
  0, 0,
  0.7579346, _,
  0, 0,
  0.7574463, _,
  0, 0,
  0.7572021, _,
  0, 0,
  0.7617188, _,
  0, 0,
  0.9388428, _,
  0, 0,
  0.9299927, _,
  0, 0,
  0.8949585, _,
  0, 0,
  0.869812, _,
  0, 0,
  0.8510132, _,
  0, 0,
  0.8327637, _,
  0, 0,
  0.8169556, _,
  0, 0,
  0.8040771, _,
  0, 0,
  0.793396, _,
  0, 0,
  0.7841797, _,
  0, 0,
  0.7803345, _,
  0, 0,
  0.7817993, _,
  0, 0,
  0.7821655, _,
  0, 0,
  0.7783203, _,
  0, 0,
  0.774231, _,
  0, 0,
  0.8469238, _,
  0, 0,
  1.046631, _,
  0, 0,
  1.005371, _,
  0, 0,
  0.975769, _,
  0, 0,
  0.9517212, _,
  0, 0,
  0.9257812, _,
  0, 0,
  0.9033813, _,
  0, 0,
  1.107117, _,
  0, 0,
  1.307861, _,
  0, 0,
  1.261475, _,
  0, 0,
  1.257568, _,
  0, 0,
  1.222717, _,
  0, 0,
  1.335938, _,
  0, 0,
  1.45874, _,
  0, 0,
  1.444275, _,
  0, 0,
  1.408447, _,
  0, 0,
  1.506287, _,
  0, 0,
  1.521118, _,
  0, 0,
  1.484802, _,
  0, 0,
  1.431335, _,
  0, 0,
  1.559998, _,
  0, 0,
  1.657654, _,
  0, 0,
  2.927979, _,
  0, 0,
  2.836792, _,
  0, 0,
  2.718567, _,
  0, 0,
  2.627197, _,
  0, 0,
  2.495911, _,
  0, 0,
  2.369263, _,
  0, 0,
  2.892639, _,
  0, 0,
  3.645569, _,
  0, 0,
  10.22552, _,
  0, 0,
  12.07367, _,
  0, 0,
  12.32074, _,
  0, 0,
  14.27448, _,
  0, 0,
  15.7373, _,
  0, 0,
  15.62836, _,
  0, 0,
  14.8349, _,
  0, 0,
  14.21692, _,
  0, 0,
  13.49945, _,
  0, 0,
  14.35162, _,
  0, 0,
  13.8584, _,
  0, 0,
  13.76477, _,
  0, 0,
  13.9303, _,
  0, 0,
  12.99426, _,
  0, 0,
  12.74249, _,
  0, 0,
  16.9043, _,
  0, 0,
  16.66034, _,
  0, 0,
  16.54449, _,
  0, 0,
  16.28705, _,
  0, 0,
  15.3869, _,
  0, 0,
  14.6358, _,
  0, 0,
  14.96265, _,
  0, 0,
  14.50903, _,
  0, 0,
  15.72174, _,
  0, 0,
  17.06964, _,
  0, 0,
  16.2655, _,
  0, 0,
  22.79614, _,
  0, 0,
  25.00195, _,
  0, 0,
  22.9455, _,
  0, 0,
  21.88794, _,
  0, 0,
  21.77808, _,
  0, 0,
  22.1709, _,
  0, 0,
  22.36523, _,
  0, 0,
  21.79462, _,
  0, 0,
  20.88177, _,
  0, 0,
  20.80518, _,
  0, 0,
  20.24469, _,
  0, 0,
  19.70709, _,
  0, 0,
  19.10138, _,
  0, 0,
  18.21436, _,
  0, 0,
  17.39166, _,
  0, 0,
  17.85101, _,
  0, 0,
  17.62146, _,
  0, 0,
  17.45673, _,
  0, 0,
  16.94922, _,
  0, 0,
  16.36475, _,
  0, 0,
  15.79761, _,
  0, 0,
  15.25989, _,
  0, 0,
  14.90814, _,
  0, 0,
  14.53937, _,
  0, 0,
  14.16614, _,
  0, 0,
  14.0014, _,
  0, 0,
  13.711, _,
  0, 0,
  13.23206, _,
  0, 0,
  12.62329, _,
  0, 0,
  12.7085, _,
  0, 0,
  12.60486, _,
  0, 0,
  15.1969, _,
  0, 0,
  23.06946, _,
  0, 0,
  24.12457, _,
  0, 0,
  25.39252, _,
  0, 0,
  23.25311, _,
  0, 0,
  22.33856, _,
  0, 0,
  21.63226, _,
  0, 0,
  21.02911, _,
  0, 0,
  20.37506, _,
  0, 0,
  20.58264, _,
  0, 0,
  20.90997, _,
  0, 0,
  20.41473, _,
  0, 0,
  19.81982, _,
  0, 0,
  19.40283, _,
  0, 0,
  19.09363, _,
  0, 0,
  19.70813, _,
  0, 0,
  19.50818, _,
  0, 0,
  19.13751, _,
  0, 0,
  18.91534, _,
  0, 0,
  18.52698, _,
  0, 0,
  18.1308, _,
  0, 0,
  17.69635, _,
  0, 0,
  17.12225, _,
  0, 0,
  16.61475, _,
  0, 0,
  16.48425, _,
  0, 0,
  18.73071, _,
  0, 0,
  19.0202, _,
  0, 0,
  18.41095, _,
  0, 0,
  18.02576, _,
  0, 0,
  17.70221, _,
  0, 0,
  17.29309, _,
  0, 0,
  16.88745, _,
  0, 0,
  16.09607, _,
  0, 0,
  15.47266, _,
  0, 0,
  14.48047, _,
  0, 0,
  13.55487, _,
  0, 0,
  12.90576, _,
  0, 0,
  12.23346, _,
  0, 0,
  12.78131, _,
  0, 0,
  12.8009, _,
  0, 0,
  12.37225, _,
  0, 0,
  11.98376, _,
  0, 0,
  11.64105, _,
  0, 0,
  11.27069, _,
  0, 0,
  10.7486, _,
  0, 0,
  10.20667, _,
  0, 0,
  9.619629, _,
  0, 0,
  8.935486, _,
  0, 0,
  8.311157, _,
  0, 0,
  7.761353, _,
  0, 0,
  7.266846, _,
  0, 0,
  6.958557, _,
  0, 0,
  7.053528, _,
  0, 0,
  6.957947, _,
  0, 0,
  6.826233, _,
  0, 0,
  6.89978, _,
  0, 0,
  6.71991, _,
  0, 0,
  6.844543, _,
  0, 0,
  8.143555, _,
  0, 0,
  11.10248, _,
  0, 0,
  11.4472, _,
  0, 0,
  11.20044, _,
  0, 0,
  12.12506, _,
  0, 0,
  26.43408, _,
  0, 0,
  26.21143, _,
  0, 0,
  26.94202, _,
  0, 0,
  25.40674, _,
  0, 0,
  23.8924, _,
  0, 0,
  22.71857, _,
  0, 0,
  21.76624, _,
  0, 0,
  21.37134, _,
  0, 0,
  20.91974, _,
  0, 0,
  20.02344, _,
  0, 0,
  19.16205, _,
  0, 0,
  19.00305, _,
  0, 0,
  18.99896, _,
  0, 0,
  17.91589, _,
  0, 0,
  16.91974, _,
  0, 0,
  15.93951, _,
  0, 0,
  14.89105, _,
  0, 0,
  13.86566, _,
  0, 0,
  12.72614, _,
  0, 0,
  13.42261, _,
  0, 0,
  21.25299, _,
  0, 0,
  22.3902, _,
  0, 0,
  21.01758, _,
  0, 0,
  19.62585, _,
  0, 0,
  18.37842, _,
  0, 0,
  17.13519, _,
  0, 0,
  15.87335, _,
  0, 0,
  14.62195, _,
  0, 0,
  13.42303, _,
  0, 0,
  12.39447, _,
  0, 0,
  11.43695, _,
  0, 0,
  11.11121, _,
  0, 0,
  10.38184, _,
  0, 0,
  9.428406, _,
  0, 0,
  8.669189, _,
  0, 0,
  7.809082, _,
  0, 0,
  6.823547, _,
  0, 0,
  6.06427, _,
  0, 0,
  5.560303, _,
  0, 0,
  5.150574, _,
  0, 0,
  4.728821, _,
  0, 0,
  4.34259, _,
  0, 0,
  4.048706, _,
  0, 0,
  3.760437, _,
  0, 0,
  3.632141, _,
  0, 0,
  3.5495, _,
  0, 0,
  3.538818, _,
  0, 0,
  4.102051, _,
  0, 0,
  4.290222, _,
  0, 0,
  4.046509, _,
  0, 0,
  3.719482, _,
  0, 0,
  3.414246, _,
  0, 0,
  3.137207, _,
  0, 0,
  2.897705, _,
  0, 0,
  2.689209, _,
  0, 0,
  2.513184, _,
  0, 0,
  2.51532, _,
  0, 0,
  2.723511, _,
  0, 0,
  2.722656, _,
  0, 0,
  2.58551, _,
  0, 0,
  2.414001, _,
  0, 0,
  2.642944, _,
  0, 0,
  4.217163, _,
  0, 0,
  4.551086, _,
  0, 0,
  5.098022, _,
  0, 0,
  6.303711, _,
  0, 0,
  6.115967, _,
  0, 0,
  5.647095, _,
  0, 0,
  5.911255, _,
  0, 0,
  6.323669, _,
  0, 0,
  6.768066, _,
  0, 0,
  6.736816, _,
  0, 0,
  6.749939, _,
  0, 0,
  6.032837, _,
  0, 0,
  5.844543, _,
  0, 0,
  5.681641, _,
  0, 0,
  7.834717, _,
  0, 0,
  11.43469, _,
  0, 0,
  10.11633, _,
  0, 0,
  9.02533, _,
  0, 0,
  7.657104, _,
  0, 0,
  17.34766, _,
  0, 0,
  24.31409, _,
  0, 0,
  28.66626, _,
  0, 0,
  26.18958, _,
  0, 0,
  23.47571, _,
  0, 0,
  21.02997, _,
  0, 0,
  18.883, _,
  0, 0,
  17.38312, _,
  0, 0,
  15.53186, _,
  0, 0,
  13.37085, _,
  0, 0,
  11.45026, _,
  0, 0,
  10.70667, _,
  0, 0,
  10.17438, _,
  0, 0,
  9.81604, _,
  0, 0,
  13.11499, _,
  0, 0,
  11.69287, _,
  0, 0,
  9.900085, _,
  0, 0,
  10.30579, _,
  0, 0,
  16.83154, _,
  0, 0,
  25.6969, _,
  0, 0,
  29.92963, _,
  0, 0,
  27.0343, _,
  0, 0,
  24.95093, _,
  0, 0,
  22.74902, _,
  0, 0,
  20.55286, _,
  0, 0,
  18.10529, _,
  0, 0,
  15.07568, _,
  0, 0,
  11.85132, _,
  0, 0,
  9.087646, _,
  0, 0,
  10.66614, _,
  0, 0,
  20.7655, _,
  0, 0,
  21.39441, _,
  0, 0,
  18.45868, _,
  0, 0,
  15.52869, _,
  0, 0,
  12.89716, _,
  0, 0,
  10.87506, _,
  0, 0,
  10.21204, _,
  0, 0,
  8.683228, _,
  0, 0,
  7.003479, _,
  0, 0,
  5.541565, _,
  0, 0,
  4.648376, _,
  0, 0,
  4.90332, _,
  0, 0,
  4.701355, _,
  0, 0,
  4.163086, _,
  0, 0,
  3.557007, _,
  0, 0,
  3.096252, _,
  0, 0,
  2.808777, _,
  0, 0,
  3.594116, _,
  0, 0,
  4.677856, _,
  0, 0,
  3.971375, _,
  0, 0,
  3.378479, _,
  0, 0,
  2.938721, _,
  0, 0,
  2.671448, _,
  0, 0,
  2.629333, _,
  0, 0,
  2.998779, _,
  0, 0,
  4.594055, _,
  0, 0,
  5.625061, _,
  0, 0,
  5.885498, _,
  0, 0,
  5.685181, _,
  0, 0,
  5.621643, _,
  0, 0,
  5.098694, _,
  0, 0,
  5.118347, _,
  0, 0,
  4.374817, _,
  0, 0,
  3.58197, _,
  0, 0,
  2.975159, _,
  0, 0,
  2.528198, _,
  0, 0,
  2.233398, _,
  0, 0,
  2.048584, _,
  0, 0,
  1.922485, _,
  0, 0,
  1.846436, _,
  0, 0,
  1.781921, _,
  0, 0,
  1.714966, _,
  0, 0,
  1.671936, _,
  0, 0,
  1.625244, _,
  0, 0,
  1.583557, _,
  0, 0,
  1.563171, _,
  0, 0,
  1.560852, _,
  0, 0,
  1.564941, _,
  0, 0,
  1.561951, _,
  0, 0,
  1.547607, _,
  0, 0,
  1.529663, _,
  0, 0,
  1.503845, _,
  0, 0,
  1.47229, _,
  0, 0,
  1.442017, _,
  0, 0,
  1.458191, _,
  0, 0,
  1.608521, _,
  0, 0,
  1.562378, _,
  0, 0,
  1.469971, _,
  0, 0,
  1.420288, _,
  0, 0,
  1.3927, _,
  0, 0,
  1.368286, _,
  0, 0,
  1.35553, _,
  0, 0,
  1.356995, _,
  0, 0,
  1.368103, _,
  0, 0,
  1.356445, _,
  0, 0,
  1.344299, _,
  0, 0,
  1.327087, _,
  0, 0,
  1.305237, _,
  0, 0,
  1.285583, _,
  0, 0,
  1.272156, _,
  0, 0,
  1.261902, _,
  0, 0,
  1.248657, _,
  0, 0,
  1.228271, _,
  0, 0,
  1.214539, _,
  0, 0,
  1.229675, _,
  0, 0,
  1.23291, _,
  0, 0,
  1.219849, _,
  0, 0,
  1.255615, _,
  0, 0,
  1.249817, _,
  0, 0,
  1.236755, _,
  0, 0,
  1.233459, _,
  0, 0,
  1.237488, _,
  0, 0,
  1.851562, _,
  0, 0,
  6.73645, _,
  0, 0,
  7.96759, _,
  0, 0,
  6.668274, _,
  0, 0,
  5.41156, _,
  0, 0,
  4.463745, _,
  0, 0,
  3.736328, _,
  0, 0,
  3.186951, _,
  0, 0,
  2.769409, _,
  0, 0,
  2.430542, _,
  0, 0,
  2.158386, _,
  0, 0,
  1.989502, _,
  0, 0,
  1.89624, _,
  0, 0,
  2.052429, _,
  0, 0,
  2.157959, _,
  0, 0,
  2.298889, _,
  0, 0,
  2.199951, _,
  0, 0,
  2.054077, _,
  0, 0,
  1.923096, _,
  0, 0,
  1.858093, _,
  0, 0,
  1.987305, _,
  0, 0,
  2.000854, _,
  0, 0,
  1.899902, _,
  0, 0,
  1.776978, _,
  0, 0,
  1.660522, _,
  0, 0,
  1.568237, _,
  0, 0,
  1.502258, _,
  0, 0,
  1.451355, _,
  0, 0,
  1.402954, _,
  0, 0,
  1.375671, _,
  0, 0,
  1.429077, _,
  0, 0,
  1.532043, _,
  0, 0,
  1.604187, _,
  0, 0,
  1.619385, _,
  0, 0,
  1.619873, _,
  0, 0,
  1.583435, _,
  0, 0,
  1.526672, _,
  0, 0,
  1.467773, _,
  0, 0,
  1.416077, _,
  0, 0,
  1.398865, _,
  0, 0,
  1.494873, _,
  0, 0,
  1.56366, _,
  0, 0,
  1.50116, _,
  0, 0,
  1.434631, _,
  0, 0,
  1.382507, _,
  0, 0,
  1.333252, _,
  0, 0,
  1.344971, _,
  0, 0,
  1.326477, _,
  0, 0,
  1.286987, _,
  0, 0,
  1.253296, _,
  0, 0,
  1.262329, _,
  0, 0,
  1.475586, _,
  0, 0,
  1.822693, _,
  0, 0,
  2.601135, _,
  0, 0,
  2.457886, _,
  0, 0,
  2.318726, _,
  0, 0,
  2.196472, _,
  0, 0,
  3.103394, _,
  0, 0,
  6.408142, _,
  0, 0,
  9.246216, _,
  0, 0,
  10.41229, _,
  0, 0,
  10.12787, _,
  0, 0,
  9.578491, _,
  0, 0,
  8.880859, _,
  0, 0,
  8.193726, _,
  0, 0,
  8.12323, _,
  0, 0,
  11.85632, _,
  0, 0,
  13.09253, _,
  0, 0,
  12.62396, _,
  0, 0,
  15.17847, _,
  0, 0,
  17.01868, _,
  0, 0,
  16.0708, _,
  0, 0,
  15.6629, _,
  0, 0,
  14.78735, _,
  0, 0,
  13.98889, _,
  0, 0,
  13.4541, _,
  0, 0,
  13.216, _,
  0, 0,
  12.95709, _,
  0, 0,
  12.85992, _,
  0, 0,
  12.17926, _,
  0, 0,
  11.67535, _,
  0, 0,
  11.25085, _,
  0, 0,
  10.98627, _,
  0, 0,
  10.73999, _,
  0, 0,
  10.33752, _,
  0, 0,
  9.884155, _,
  0, 0,
  11.1214, _,
  0, 0,
  18.29272, _,
  0, 0,
  20.51819, _,
  0, 0,
  19.34497, _,
  0, 0,
  18.29669, _,
  0, 0,
  17.41925, _,
  0, 0,
  16.71552, _,
  0, 0,
  16.3689, _,
  0, 0,
  17.3894, _,
  0, 0,
  18.08826, _,
  0, 0,
  18.6261, _ ;

 time = 50400.5, 50401.5, 50402.5, 50403.5, 50404.5, 50405.5, 50406.5, 
    50407.5, 50408.5, 50409.5, 50410.5, 50411.5, 50412.5, 50413.5, 50414.5, 
    50415.5, 50416.5, 50417.5, 50418.5, 50419.5, 50420.5, 50421.5, 50422.5, 
    50423.5, 50424.5, 50425.5, 50426.5, 50427.5, 50428.5, 50429.5, 50430.5, 
    50431.5, 50432.5, 50433.5, 50434.5, 50435.5, 50436.5, 50437.5, 50438.5, 
    50439.5, 50440.5, 50441.5, 50442.5, 50443.5, 50444.5, 50445.5, 50446.5, 
    50447.5, 50448.5, 50449.5, 50450.5, 50451.5, 50452.5, 50453.5, 50454.5, 
    50455.5, 50456.5, 50457.5, 50458.5, 50459.5, 50460.5, 50461.5, 50462.5, 
    50463.5, 50464.5, 50465.5, 50466.5, 50467.5, 50468.5, 50469.5, 50470.5, 
    50471.5, 50472.5, 50473.5, 50474.5, 50475.5, 50476.5, 50477.5, 50478.5, 
    50479.5, 50480.5, 50481.5, 50482.5, 50483.5, 50484.5, 50485.5, 50486.5, 
    50487.5, 50488.5, 50489.5, 50490.5, 50491.5, 50492.5, 50493.5, 50494.5, 
    50495.5, 50496.5, 50497.5, 50498.5, 50499.5, 50500.5, 50501.5, 50502.5, 
    50503.5, 50504.5, 50505.5, 50506.5, 50507.5, 50508.5, 50509.5, 50510.5, 
    50511.5, 50512.5, 50513.5, 50514.5, 50515.5, 50516.5, 50517.5, 50518.5, 
    50519.5, 50520.5, 50521.5, 50522.5, 50523.5, 50524.5, 50525.5, 50526.5, 
    50527.5, 50528.5, 50529.5, 50530.5, 50531.5, 50532.5, 50533.5, 50534.5, 
    50535.5, 50536.5, 50537.5, 50538.5, 50539.5, 50540.5, 50541.5, 50542.5, 
    50543.5, 50544.5, 50545.5, 50546.5, 50547.5, 50548.5, 50549.5, 50550.5, 
    50551.5, 50552.5, 50553.5, 50554.5, 50555.5, 50556.5, 50557.5, 50558.5, 
    50559.5, 50560.5, 50561.5, 50562.5, 50563.5, 50564.5, 50565.5, 50566.5, 
    50567.5, 50568.5, 50569.5, 50570.5, 50571.5, 50572.5, 50573.5, 50574.5, 
    50575.5, 50576.5, 50577.5, 50578.5, 50579.5, 50580.5, 50581.5, 50582.5, 
    50583.5, 50584.5, 50585.5, 50586.5, 50587.5, 50588.5, 50589.5, 50590.5, 
    50591.5, 50592.5, 50593.5, 50594.5, 50595.5, 50596.5, 50597.5, 50598.5, 
    50599.5, 50600.5, 50601.5, 50602.5, 50603.5, 50604.5, 50605.5, 50606.5, 
    50607.5, 50608.5, 50609.5, 50610.5, 50611.5, 50612.5, 50613.5, 50614.5, 
    50615.5, 50616.5, 50617.5, 50618.5, 50619.5, 50620.5, 50621.5, 50622.5, 
    50623.5, 50624.5, 50625.5, 50626.5, 50627.5, 50628.5, 50629.5, 50630.5, 
    50631.5, 50632.5, 50633.5, 50634.5, 50635.5, 50636.5, 50637.5, 50638.5, 
    50639.5, 50640.5, 50641.5, 50642.5, 50643.5, 50644.5, 50645.5, 50646.5, 
    50647.5, 50648.5, 50649.5, 50650.5, 50651.5, 50652.5, 50653.5, 50654.5, 
    50655.5, 50656.5, 50657.5, 50658.5, 50659.5, 50660.5, 50661.5, 50662.5, 
    50663.5, 50664.5, 50665.5, 50666.5, 50667.5, 50668.5, 50669.5, 50670.5, 
    50671.5, 50672.5, 50673.5, 50674.5, 50675.5, 50676.5, 50677.5, 50678.5, 
    50679.5, 50680.5, 50681.5, 50682.5, 50683.5, 50684.5, 50685.5, 50686.5, 
    50687.5, 50688.5, 50689.5, 50690.5, 50691.5, 50692.5, 50693.5, 50694.5, 
    50695.5, 50696.5, 50697.5, 50698.5, 50699.5, 50700.5, 50701.5, 50702.5, 
    50703.5, 50704.5, 50705.5, 50706.5, 50707.5, 50708.5, 50709.5, 50710.5, 
    50711.5, 50712.5, 50713.5, 50714.5, 50715.5, 50716.5, 50717.5, 50718.5, 
    50719.5, 50720.5, 50721.5, 50722.5, 50723.5, 50724.5, 50725.5, 50726.5, 
    50727.5, 50728.5, 50729.5, 50730.5, 50731.5, 50732.5, 50733.5, 50734.5, 
    50735.5, 50736.5, 50737.5, 50738.5, 50739.5, 50740.5, 50741.5, 50742.5, 
    50743.5, 50744.5, 50745.5, 50746.5, 50747.5, 50748.5, 50749.5, 50750.5, 
    50751.5, 50752.5, 50753.5, 50754.5, 50755.5, 50756.5, 50757.5, 50758.5, 
    50759.5, 50760.5, 50761.5, 50762.5, 50763.5, 50764.5, 50765.5, 50766.5, 
    50767.5, 50768.5, 50769.5, 50770.5, 50771.5, 50772.5, 50773.5, 50774.5, 
    50775.5, 50776.5, 50777.5, 50778.5, 50779.5, 50780.5, 50781.5, 50782.5, 
    50783.5, 50784.5, 50785.5, 50786.5, 50787.5, 50788.5, 50789.5, 50790.5, 
    50791.5, 50792.5, 50793.5, 50794.5, 50795.5, 50796.5, 50797.5, 50798.5, 
    50799.5, 50800.5, 50801.5, 50802.5, 50803.5, 50804.5, 50805.5, 50806.5, 
    50807.5, 50808.5, 50809.5, 50810.5, 50811.5, 50812.5, 50813.5, 50814.5, 
    50815.5, 50816.5, 50817.5, 50818.5, 50819.5, 50820.5, 50821.5, 50822.5, 
    50823.5, 50824.5, 50825.5, 50826.5, 50827.5, 50828.5, 50829.5, 50830.5, 
    50831.5, 50832.5, 50833.5, 50834.5, 50835.5, 50836.5, 50837.5, 50838.5, 
    50839.5, 50840.5, 50841.5, 50842.5, 50843.5, 50844.5, 50845.5, 50846.5, 
    50847.5, 50848.5, 50849.5, 50850.5, 50851.5, 50852.5, 50853.5, 50854.5, 
    50855.5, 50856.5, 50857.5, 50858.5, 50859.5, 50860.5, 50861.5, 50862.5, 
    50863.5, 50864.5, 50865.5, 50866.5, 50867.5, 50868.5, 50869.5, 50870.5, 
    50871.5, 50872.5, 50873.5, 50874.5, 50875.5, 50876.5, 50877.5, 50878.5, 
    50879.5, 50880.5, 50881.5, 50882.5, 50883.5, 50884.5, 50885.5, 50886.5, 
    50887.5, 50888.5, 50889.5, 50890.5, 50891.5, 50892.5, 50893.5, 50894.5, 
    50895.5, 50896.5, 50897.5, 50898.5, 50899.5, 50900.5, 50901.5, 50902.5, 
    50903.5, 50904.5, 50905.5, 50906.5, 50907.5, 50908.5, 50909.5, 50910.5, 
    50911.5, 50912.5, 50913.5, 50914.5, 50915.5, 50916.5, 50917.5, 50918.5, 
    50919.5, 50920.5, 50921.5, 50922.5, 50923.5, 50924.5, 50925.5, 50926.5, 
    50927.5, 50928.5, 50929.5, 50930.5, 50931.5, 50932.5, 50933.5, 50934.5, 
    50935.5, 50936.5, 50937.5, 50938.5, 50939.5, 50940.5, 50941.5, 50942.5, 
    50943.5, 50944.5, 50945.5, 50946.5, 50947.5, 50948.5, 50949.5, 50950.5, 
    50951.5, 50952.5, 50953.5, 50954.5, 50955.5, 50956.5, 50957.5, 50958.5, 
    50959.5, 50960.5, 50961.5, 50962.5, 50963.5, 50964.5, 50965.5, 50966.5, 
    50967.5, 50968.5, 50969.5, 50970.5, 50971.5, 50972.5, 50973.5, 50974.5, 
    50975.5, 50976.5, 50977.5, 50978.5, 50979.5, 50980.5, 50981.5, 50982.5, 
    50983.5, 50984.5, 50985.5, 50986.5, 50987.5, 50988.5, 50989.5, 50990.5, 
    50991.5, 50992.5, 50993.5, 50994.5, 50995.5, 50996.5, 50997.5, 50998.5, 
    50999.5, 51000.5, 51001.5, 51002.5, 51003.5, 51004.5, 51005.5, 51006.5, 
    51007.5, 51008.5, 51009.5, 51010.5, 51011.5, 51012.5, 51013.5, 51014.5, 
    51015.5, 51016.5, 51017.5, 51018.5, 51019.5, 51020.5, 51021.5, 51022.5, 
    51023.5, 51024.5, 51025.5, 51026.5, 51027.5, 51028.5, 51029.5, 51030.5, 
    51031.5, 51032.5, 51033.5, 51034.5, 51035.5, 51036.5, 51037.5, 51038.5, 
    51039.5, 51040.5, 51041.5, 51042.5, 51043.5, 51044.5, 51045.5, 51046.5, 
    51047.5, 51048.5, 51049.5, 51050.5, 51051.5, 51052.5, 51053.5, 51054.5, 
    51055.5, 51056.5, 51057.5, 51058.5, 51059.5, 51060.5, 51061.5, 51062.5, 
    51063.5, 51064.5, 51065.5, 51066.5, 51067.5, 51068.5, 51069.5, 51070.5, 
    51071.5, 51072.5, 51073.5, 51074.5, 51075.5, 51076.5, 51077.5, 51078.5, 
    51079.5, 51080.5, 51081.5, 51082.5, 51083.5, 51084.5, 51085.5, 51086.5, 
    51087.5, 51088.5, 51089.5, 51090.5, 51091.5, 51092.5, 51093.5, 51094.5, 
    51095.5, 51096.5, 51097.5, 51098.5, 51099.5, 51100.5, 51101.5, 51102.5, 
    51103.5, 51104.5, 51105.5, 51106.5, 51107.5, 51108.5, 51109.5, 51110.5, 
    51111.5, 51112.5, 51113.5, 51114.5, 51115.5, 51116.5, 51117.5, 51118.5, 
    51119.5, 51120.5, 51121.5, 51122.5, 51123.5, 51124.5, 51125.5, 51126.5, 
    51127.5, 51128.5, 51129.5, 51130.5, 51131.5, 51132.5, 51133.5, 51134.5, 
    51135.5, 51136.5, 51137.5, 51138.5, 51139.5, 51140.5, 51141.5, 51142.5, 
    51143.5, 51144.5, 51145.5, 51146.5, 51147.5, 51148.5, 51149.5, 51150.5, 
    51151.5, 51152.5, 51153.5, 51154.5, 51155.5, 51156.5, 51157.5, 51158.5, 
    51159.5, 51160.5, 51161.5, 51162.5, 51163.5, 51164.5, 51165.5, 51166.5, 
    51167.5, 51168.5, 51169.5, 51170.5, 51171.5, 51172.5, 51173.5, 51174.5, 
    51175.5, 51176.5, 51177.5, 51178.5, 51179.5, 51180.5, 51181.5, 51182.5, 
    51183.5, 51184.5, 51185.5, 51186.5, 51187.5, 51188.5, 51189.5, 51190.5, 
    51191.5, 51192.5, 51193.5, 51194.5, 51195.5, 51196.5, 51197.5, 51198.5, 
    51199.5, 51200.5, 51201.5, 51202.5, 51203.5, 51204.5, 51205.5, 51206.5, 
    51207.5, 51208.5, 51209.5, 51210.5, 51211.5, 51212.5, 51213.5, 51214.5, 
    51215.5, 51216.5, 51217.5, 51218.5, 51219.5, 51220.5, 51221.5, 51222.5, 
    51223.5, 51224.5, 51225.5, 51226.5, 51227.5, 51228.5, 51229.5, 51230.5, 
    51231.5, 51232.5, 51233.5, 51234.5, 51235.5, 51236.5, 51237.5, 51238.5, 
    51239.5, 51240.5, 51241.5, 51242.5, 51243.5, 51244.5, 51245.5, 51246.5, 
    51247.5, 51248.5, 51249.5, 51250.5, 51251.5, 51252.5, 51253.5, 51254.5, 
    51255.5, 51256.5, 51257.5, 51258.5, 51259.5, 51260.5, 51261.5, 51262.5, 
    51263.5, 51264.5, 51265.5, 51266.5, 51267.5, 51268.5, 51269.5, 51270.5, 
    51271.5, 51272.5, 51273.5, 51274.5, 51275.5, 51276.5, 51277.5, 51278.5, 
    51279.5, 51280.5, 51281.5, 51282.5, 51283.5, 51284.5, 51285.5, 51286.5, 
    51287.5, 51288.5, 51289.5, 51290.5, 51291.5, 51292.5, 51293.5, 51294.5, 
    51295.5, 51296.5, 51297.5, 51298.5, 51299.5, 51300.5, 51301.5, 51302.5, 
    51303.5, 51304.5, 51305.5, 51306.5, 51307.5, 51308.5, 51309.5, 51310.5, 
    51311.5, 51312.5, 51313.5, 51314.5, 51315.5, 51316.5, 51317.5, 51318.5, 
    51319.5, 51320.5, 51321.5, 51322.5, 51323.5, 51324.5, 51325.5, 51326.5, 
    51327.5, 51328.5, 51329.5, 51330.5, 51331.5, 51332.5, 51333.5, 51334.5, 
    51335.5, 51336.5, 51337.5, 51338.5, 51339.5, 51340.5, 51341.5, 51342.5, 
    51343.5, 51344.5, 51345.5, 51346.5, 51347.5, 51348.5, 51349.5, 51350.5, 
    51351.5, 51352.5, 51353.5, 51354.5, 51355.5, 51356.5, 51357.5, 51358.5, 
    51359.5, 51360.5, 51361.5, 51362.5, 51363.5, 51364.5, 51365.5, 51366.5, 
    51367.5, 51368.5, 51369.5, 51370.5, 51371.5, 51372.5, 51373.5, 51374.5, 
    51375.5, 51376.5, 51377.5, 51378.5, 51379.5, 51380.5, 51381.5, 51382.5, 
    51383.5, 51384.5, 51385.5, 51386.5, 51387.5, 51388.5, 51389.5, 51390.5, 
    51391.5, 51392.5, 51393.5, 51394.5, 51395.5, 51396.5, 51397.5, 51398.5, 
    51399.5, 51400.5, 51401.5, 51402.5, 51403.5, 51404.5, 51405.5, 51406.5, 
    51407.5, 51408.5, 51409.5, 51410.5, 51411.5, 51412.5, 51413.5, 51414.5, 
    51415.5, 51416.5, 51417.5, 51418.5, 51419.5, 51420.5, 51421.5, 51422.5, 
    51423.5, 51424.5, 51425.5, 51426.5, 51427.5, 51428.5, 51429.5, 51430.5, 
    51431.5, 51432.5, 51433.5, 51434.5, 51435.5, 51436.5, 51437.5, 51438.5, 
    51439.5, 51440.5, 51441.5, 51442.5, 51443.5, 51444.5, 51445.5, 51446.5, 
    51447.5, 51448.5, 51449.5, 51450.5, 51451.5, 51452.5, 51453.5, 51454.5, 
    51455.5, 51456.5, 51457.5, 51458.5, 51459.5, 51460.5, 51461.5, 51462.5, 
    51463.5, 51464.5, 51465.5, 51466.5, 51467.5, 51468.5, 51469.5, 51470.5, 
    51471.5, 51472.5, 51473.5, 51474.5, 51475.5, 51476.5, 51477.5, 51478.5, 
    51479.5, 51480.5, 51481.5, 51482.5, 51483.5, 51484.5, 51485.5, 51486.5, 
    51487.5, 51488.5, 51489.5, 51490.5, 51491.5, 51492.5, 51493.5, 51494.5, 
    51495.5, 51496.5, 51497.5, 51498.5, 51499.5, 51500.5, 51501.5, 51502.5, 
    51503.5, 51504.5, 51505.5, 51506.5, 51507.5, 51508.5, 51509.5, 51510.5, 
    51511.5, 51512.5, 51513.5, 51514.5, 51515.5, 51516.5, 51517.5, 51518.5, 
    51519.5, 51520.5, 51521.5, 51522.5, 51523.5, 51524.5, 51525.5, 51526.5, 
    51527.5, 51528.5, 51529.5, 51530.5, 51531.5, 51532.5, 51533.5, 51534.5, 
    51535.5, 51536.5, 51537.5, 51538.5, 51539.5, 51540.5, 51541.5, 51542.5, 
    51543.5, 51544.5, 51545.5, 51546.5, 51547.5, 51548.5, 51549.5, 51550.5, 
    51551.5, 51552.5, 51553.5, 51554.5, 51555.5, 51556.5, 51557.5, 51558.5, 
    51559.5, 51560.5, 51561.5, 51562.5, 51563.5, 51564.5, 51565.5, 51566.5, 
    51567.5, 51568.5, 51569.5, 51570.5, 51571.5, 51572.5, 51573.5, 51574.5, 
    51575.5, 51576.5, 51577.5, 51578.5, 51579.5, 51580.5, 51581.5, 51582.5, 
    51583.5, 51584.5, 51585.5, 51586.5, 51587.5, 51588.5, 51589.5, 51590.5, 
    51591.5, 51592.5, 51593.5, 51594.5, 51595.5, 51596.5, 51597.5, 51598.5, 
    51599.5, 51600.5, 51601.5, 51602.5, 51603.5, 51604.5, 51605.5, 51606.5, 
    51607.5, 51608.5, 51609.5, 51610.5, 51611.5, 51612.5, 51613.5, 51614.5, 
    51615.5, 51616.5, 51617.5, 51618.5, 51619.5, 51620.5, 51621.5, 51622.5, 
    51623.5, 51624.5, 51625.5, 51626.5, 51627.5, 51628.5, 51629.5, 51630.5, 
    51631.5, 51632.5, 51633.5, 51634.5, 51635.5, 51636.5, 51637.5, 51638.5, 
    51639.5, 51640.5, 51641.5, 51642.5, 51643.5, 51644.5, 51645.5, 51646.5, 
    51647.5, 51648.5, 51649.5, 51650.5, 51651.5, 51652.5, 51653.5, 51654.5, 
    51655.5, 51656.5, 51657.5, 51658.5, 51659.5, 51660.5, 51661.5, 51662.5, 
    51663.5, 51664.5, 51665.5, 51666.5, 51667.5, 51668.5, 51669.5, 51670.5, 
    51671.5, 51672.5, 51673.5, 51674.5, 51675.5, 51676.5, 51677.5, 51678.5, 
    51679.5, 51680.5, 51681.5, 51682.5, 51683.5, 51684.5, 51685.5, 51686.5, 
    51687.5, 51688.5, 51689.5, 51690.5, 51691.5, 51692.5, 51693.5, 51694.5, 
    51695.5, 51696.5, 51697.5, 51698.5, 51699.5, 51700.5, 51701.5, 51702.5, 
    51703.5, 51704.5, 51705.5, 51706.5, 51707.5, 51708.5, 51709.5, 51710.5, 
    51711.5, 51712.5, 51713.5, 51714.5, 51715.5, 51716.5, 51717.5, 51718.5, 
    51719.5, 51720.5, 51721.5, 51722.5, 51723.5, 51724.5, 51725.5, 51726.5, 
    51727.5, 51728.5, 51729.5, 51730.5, 51731.5, 51732.5, 51733.5, 51734.5, 
    51735.5, 51736.5, 51737.5, 51738.5, 51739.5, 51740.5, 51741.5, 51742.5, 
    51743.5, 51744.5, 51745.5, 51746.5, 51747.5, 51748.5, 51749.5, 51750.5, 
    51751.5, 51752.5, 51753.5, 51754.5, 51755.5, 51756.5, 51757.5, 51758.5, 
    51759.5, 51760.5, 51761.5, 51762.5, 51763.5, 51764.5, 51765.5, 51766.5, 
    51767.5, 51768.5, 51769.5, 51770.5, 51771.5, 51772.5, 51773.5, 51774.5, 
    51775.5, 51776.5, 51777.5, 51778.5, 51779.5, 51780.5, 51781.5, 51782.5, 
    51783.5, 51784.5, 51785.5, 51786.5, 51787.5, 51788.5, 51789.5, 51790.5, 
    51791.5, 51792.5, 51793.5, 51794.5, 51795.5, 51796.5, 51797.5, 51798.5, 
    51799.5, 51800.5, 51801.5, 51802.5, 51803.5, 51804.5, 51805.5, 51806.5, 
    51807.5, 51808.5, 51809.5, 51810.5, 51811.5, 51812.5, 51813.5, 51814.5, 
    51815.5, 51816.5, 51817.5, 51818.5, 51819.5, 51820.5, 51821.5, 51822.5, 
    51823.5, 51824.5, 51825.5, 51826.5, 51827.5, 51828.5, 51829.5, 51830.5, 
    51831.5, 51832.5, 51833.5, 51834.5, 51835.5, 51836.5, 51837.5, 51838.5, 
    51839.5, 51840.5, 51841.5, 51842.5, 51843.5, 51844.5, 51845.5, 51846.5, 
    51847.5, 51848.5, 51849.5, 51850.5, 51851.5, 51852.5, 51853.5, 51854.5, 
    51855.5, 51856.5, 51857.5, 51858.5, 51859.5, 51860.5, 51861.5, 51862.5, 
    51863.5, 51864.5, 51865.5, 51866.5, 51867.5, 51868.5, 51869.5, 51870.5, 
    51871.5, 51872.5, 51873.5, 51874.5, 51875.5, 51876.5, 51877.5, 51878.5, 
    51879.5, 51880.5, 51881.5, 51882.5, 51883.5, 51884.5, 51885.5, 51886.5, 
    51887.5, 51888.5, 51889.5, 51890.5, 51891.5, 51892.5, 51893.5, 51894.5, 
    51895.5, 51896.5, 51897.5, 51898.5, 51899.5, 51900.5, 51901.5, 51902.5, 
    51903.5, 51904.5, 51905.5, 51906.5, 51907.5, 51908.5, 51909.5, 51910.5, 
    51911.5, 51912.5, 51913.5, 51914.5, 51915.5, 51916.5, 51917.5, 51918.5, 
    51919.5, 51920.5, 51921.5, 51922.5, 51923.5, 51924.5, 51925.5, 51926.5, 
    51927.5, 51928.5, 51929.5, 51930.5, 51931.5, 51932.5, 51933.5, 51934.5, 
    51935.5, 51936.5, 51937.5, 51938.5, 51939.5, 51940.5, 51941.5, 51942.5, 
    51943.5, 51944.5, 51945.5, 51946.5, 51947.5, 51948.5, 51949.5, 51950.5, 
    51951.5, 51952.5, 51953.5, 51954.5, 51955.5, 51956.5, 51957.5, 51958.5, 
    51959.5, 51960.5, 51961.5, 51962.5, 51963.5, 51964.5, 51965.5, 51966.5, 
    51967.5, 51968.5, 51969.5, 51970.5, 51971.5, 51972.5, 51973.5, 51974.5, 
    51975.5, 51976.5, 51977.5, 51978.5, 51979.5, 51980.5, 51981.5, 51982.5, 
    51983.5, 51984.5, 51985.5, 51986.5, 51987.5, 51988.5, 51989.5, 51990.5, 
    51991.5, 51992.5, 51993.5, 51994.5, 51995.5, 51996.5, 51997.5, 51998.5, 
    51999.5, 52000.5, 52001.5, 52002.5, 52003.5, 52004.5, 52005.5, 52006.5, 
    52007.5, 52008.5, 52009.5, 52010.5, 52011.5, 52012.5, 52013.5, 52014.5, 
    52015.5, 52016.5, 52017.5, 52018.5, 52019.5, 52020.5, 52021.5, 52022.5, 
    52023.5, 52024.5, 52025.5, 52026.5, 52027.5, 52028.5, 52029.5, 52030.5, 
    52031.5, 52032.5, 52033.5, 52034.5, 52035.5, 52036.5, 52037.5, 52038.5, 
    52039.5, 52040.5, 52041.5, 52042.5, 52043.5, 52044.5, 52045.5, 52046.5, 
    52047.5, 52048.5, 52049.5, 52050.5, 52051.5, 52052.5, 52053.5, 52054.5, 
    52055.5, 52056.5, 52057.5, 52058.5, 52059.5, 52060.5, 52061.5, 52062.5, 
    52063.5, 52064.5, 52065.5, 52066.5, 52067.5, 52068.5, 52069.5, 52070.5, 
    52071.5, 52072.5, 52073.5, 52074.5, 52075.5, 52076.5, 52077.5, 52078.5, 
    52079.5, 52080.5, 52081.5, 52082.5, 52083.5, 52084.5, 52085.5, 52086.5, 
    52087.5, 52088.5, 52089.5, 52090.5, 52091.5, 52092.5, 52093.5, 52094.5, 
    52095.5, 52096.5, 52097.5, 52098.5, 52099.5, 52100.5, 52101.5, 52102.5, 
    52103.5, 52104.5, 52105.5, 52106.5, 52107.5, 52108.5, 52109.5, 52110.5, 
    52111.5, 52112.5, 52113.5, 52114.5, 52115.5, 52116.5, 52117.5, 52118.5, 
    52119.5, 52120.5, 52121.5, 52122.5, 52123.5, 52124.5, 52125.5, 52126.5, 
    52127.5, 52128.5, 52129.5, 52130.5, 52131.5, 52132.5, 52133.5, 52134.5, 
    52135.5, 52136.5, 52137.5, 52138.5, 52139.5, 52140.5, 52141.5, 52142.5, 
    52143.5, 52144.5, 52145.5, 52146.5, 52147.5, 52148.5, 52149.5, 52150.5, 
    52151.5, 52152.5, 52153.5, 52154.5, 52155.5, 52156.5, 52157.5, 52158.5, 
    52159.5, 52160.5, 52161.5, 52162.5, 52163.5, 52164.5, 52165.5, 52166.5, 
    52167.5, 52168.5, 52169.5, 52170.5, 52171.5, 52172.5, 52173.5, 52174.5, 
    52175.5, 52176.5, 52177.5, 52178.5, 52179.5, 52180.5, 52181.5, 52182.5, 
    52183.5, 52184.5, 52185.5, 52186.5, 52187.5, 52188.5, 52189.5, 52190.5, 
    52191.5, 52192.5, 52193.5, 52194.5, 52195.5, 52196.5, 52197.5, 52198.5, 
    52199.5, 52200.5, 52201.5, 52202.5, 52203.5, 52204.5, 52205.5, 52206.5, 
    52207.5, 52208.5, 52209.5, 52210.5, 52211.5, 52212.5, 52213.5, 52214.5, 
    52215.5, 52216.5, 52217.5, 52218.5, 52219.5, 52220.5, 52221.5, 52222.5, 
    52223.5, 52224.5, 52225.5, 52226.5, 52227.5, 52228.5, 52229.5, 52230.5, 
    52231.5, 52232.5, 52233.5, 52234.5, 52235.5, 52236.5, 52237.5, 52238.5, 
    52239.5, 52240.5, 52241.5, 52242.5, 52243.5, 52244.5, 52245.5, 52246.5, 
    52247.5, 52248.5, 52249.5, 52250.5, 52251.5, 52252.5, 52253.5, 52254.5, 
    52255.5, 52256.5, 52257.5, 52258.5, 52259.5, 52260.5, 52261.5, 52262.5, 
    52263.5, 52264.5, 52265.5, 52266.5, 52267.5, 52268.5, 52269.5, 52270.5, 
    52271.5, 52272.5, 52273.5, 52274.5, 52275.5, 52276.5, 52277.5, 52278.5, 
    52279.5, 52280.5, 52281.5, 52282.5, 52283.5, 52284.5, 52285.5, 52286.5, 
    52287.5, 52288.5, 52289.5, 52290.5, 52291.5, 52292.5, 52293.5, 52294.5, 
    52295.5, 52296.5, 52297.5, 52298.5, 52299.5, 52300.5, 52301.5, 52302.5, 
    52303.5, 52304.5, 52305.5, 52306.5, 52307.5, 52308.5, 52309.5, 52310.5, 
    52311.5, 52312.5, 52313.5, 52314.5, 52315.5, 52316.5, 52317.5, 52318.5, 
    52319.5, 52320.5, 52321.5, 52322.5, 52323.5, 52324.5, 52325.5, 52326.5, 
    52327.5, 52328.5, 52329.5, 52330.5, 52331.5, 52332.5, 52333.5, 52334.5, 
    52335.5, 52336.5, 52337.5, 52338.5, 52339.5, 52340.5, 52341.5, 52342.5, 
    52343.5, 52344.5, 52345.5, 52346.5, 52347.5, 52348.5, 52349.5, 52350.5, 
    52351.5, 52352.5, 52353.5, 52354.5, 52355.5, 52356.5, 52357.5, 52358.5, 
    52359.5, 52360.5, 52361.5, 52362.5, 52363.5, 52364.5, 52365.5, 52366.5, 
    52367.5, 52368.5, 52369.5, 52370.5, 52371.5, 52372.5, 52373.5, 52374.5, 
    52375.5, 52376.5, 52377.5, 52378.5, 52379.5, 52380.5, 52381.5, 52382.5, 
    52383.5, 52384.5, 52385.5, 52386.5, 52387.5, 52388.5, 52389.5, 52390.5, 
    52391.5, 52392.5, 52393.5, 52394.5, 52395.5, 52396.5, 52397.5, 52398.5, 
    52399.5, 52400.5, 52401.5, 52402.5, 52403.5, 52404.5, 52405.5, 52406.5, 
    52407.5, 52408.5, 52409.5, 52410.5, 52411.5, 52412.5, 52413.5, 52414.5, 
    52415.5, 52416.5, 52417.5, 52418.5, 52419.5, 52420.5, 52421.5, 52422.5, 
    52423.5, 52424.5, 52425.5, 52426.5, 52427.5, 52428.5, 52429.5, 52430.5, 
    52431.5, 52432.5, 52433.5, 52434.5, 52435.5, 52436.5, 52437.5, 52438.5, 
    52439.5, 52440.5, 52441.5, 52442.5, 52443.5, 52444.5, 52445.5, 52446.5, 
    52447.5, 52448.5, 52449.5, 52450.5, 52451.5, 52452.5, 52453.5, 52454.5, 
    52455.5, 52456.5, 52457.5, 52458.5, 52459.5, 52460.5, 52461.5, 52462.5, 
    52463.5, 52464.5, 52465.5, 52466.5, 52467.5, 52468.5, 52469.5, 52470.5, 
    52471.5, 52472.5, 52473.5, 52474.5, 52475.5, 52476.5, 52477.5, 52478.5, 
    52479.5, 52480.5, 52481.5, 52482.5, 52483.5, 52484.5, 52485.5, 52486.5, 
    52487.5, 52488.5, 52489.5, 52490.5, 52491.5, 52492.5, 52493.5, 52494.5, 
    52495.5, 52496.5, 52497.5, 52498.5, 52499.5, 52500.5, 52501.5, 52502.5, 
    52503.5, 52504.5, 52505.5, 52506.5, 52507.5, 52508.5, 52509.5, 52510.5, 
    52511.5, 52512.5, 52513.5, 52514.5, 52515.5, 52516.5, 52517.5, 52518.5, 
    52519.5, 52520.5, 52521.5, 52522.5, 52523.5, 52524.5, 52525.5, 52526.5, 
    52527.5, 52528.5, 52529.5, 52530.5, 52531.5, 52532.5, 52533.5, 52534.5, 
    52535.5, 52536.5, 52537.5, 52538.5, 52539.5, 52540.5, 52541.5, 52542.5, 
    52543.5, 52544.5, 52545.5, 52546.5, 52547.5, 52548.5, 52549.5, 52550.5, 
    52551.5, 52552.5, 52553.5, 52554.5, 52555.5, 52556.5, 52557.5, 52558.5, 
    52559.5 ;

 time_bnds =
  50400, 50401,
  50401, 50402,
  50402, 50403,
  50403, 50404,
  50404, 50405,
  50405, 50406,
  50406, 50407,
  50407, 50408,
  50408, 50409,
  50409, 50410,
  50410, 50411,
  50411, 50412,
  50412, 50413,
  50413, 50414,
  50414, 50415,
  50415, 50416,
  50416, 50417,
  50417, 50418,
  50418, 50419,
  50419, 50420,
  50420, 50421,
  50421, 50422,
  50422, 50423,
  50423, 50424,
  50424, 50425,
  50425, 50426,
  50426, 50427,
  50427, 50428,
  50428, 50429,
  50429, 50430,
  50430, 50431,
  50431, 50432,
  50432, 50433,
  50433, 50434,
  50434, 50435,
  50435, 50436,
  50436, 50437,
  50437, 50438,
  50438, 50439,
  50439, 50440,
  50440, 50441,
  50441, 50442,
  50442, 50443,
  50443, 50444,
  50444, 50445,
  50445, 50446,
  50446, 50447,
  50447, 50448,
  50448, 50449,
  50449, 50450,
  50450, 50451,
  50451, 50452,
  50452, 50453,
  50453, 50454,
  50454, 50455,
  50455, 50456,
  50456, 50457,
  50457, 50458,
  50458, 50459,
  50459, 50460,
  50460, 50461,
  50461, 50462,
  50462, 50463,
  50463, 50464,
  50464, 50465,
  50465, 50466,
  50466, 50467,
  50467, 50468,
  50468, 50469,
  50469, 50470,
  50470, 50471,
  50471, 50472,
  50472, 50473,
  50473, 50474,
  50474, 50475,
  50475, 50476,
  50476, 50477,
  50477, 50478,
  50478, 50479,
  50479, 50480,
  50480, 50481,
  50481, 50482,
  50482, 50483,
  50483, 50484,
  50484, 50485,
  50485, 50486,
  50486, 50487,
  50487, 50488,
  50488, 50489,
  50489, 50490,
  50490, 50491,
  50491, 50492,
  50492, 50493,
  50493, 50494,
  50494, 50495,
  50495, 50496,
  50496, 50497,
  50497, 50498,
  50498, 50499,
  50499, 50500,
  50500, 50501,
  50501, 50502,
  50502, 50503,
  50503, 50504,
  50504, 50505,
  50505, 50506,
  50506, 50507,
  50507, 50508,
  50508, 50509,
  50509, 50510,
  50510, 50511,
  50511, 50512,
  50512, 50513,
  50513, 50514,
  50514, 50515,
  50515, 50516,
  50516, 50517,
  50517, 50518,
  50518, 50519,
  50519, 50520,
  50520, 50521,
  50521, 50522,
  50522, 50523,
  50523, 50524,
  50524, 50525,
  50525, 50526,
  50526, 50527,
  50527, 50528,
  50528, 50529,
  50529, 50530,
  50530, 50531,
  50531, 50532,
  50532, 50533,
  50533, 50534,
  50534, 50535,
  50535, 50536,
  50536, 50537,
  50537, 50538,
  50538, 50539,
  50539, 50540,
  50540, 50541,
  50541, 50542,
  50542, 50543,
  50543, 50544,
  50544, 50545,
  50545, 50546,
  50546, 50547,
  50547, 50548,
  50548, 50549,
  50549, 50550,
  50550, 50551,
  50551, 50552,
  50552, 50553,
  50553, 50554,
  50554, 50555,
  50555, 50556,
  50556, 50557,
  50557, 50558,
  50558, 50559,
  50559, 50560,
  50560, 50561,
  50561, 50562,
  50562, 50563,
  50563, 50564,
  50564, 50565,
  50565, 50566,
  50566, 50567,
  50567, 50568,
  50568, 50569,
  50569, 50570,
  50570, 50571,
  50571, 50572,
  50572, 50573,
  50573, 50574,
  50574, 50575,
  50575, 50576,
  50576, 50577,
  50577, 50578,
  50578, 50579,
  50579, 50580,
  50580, 50581,
  50581, 50582,
  50582, 50583,
  50583, 50584,
  50584, 50585,
  50585, 50586,
  50586, 50587,
  50587, 50588,
  50588, 50589,
  50589, 50590,
  50590, 50591,
  50591, 50592,
  50592, 50593,
  50593, 50594,
  50594, 50595,
  50595, 50596,
  50596, 50597,
  50597, 50598,
  50598, 50599,
  50599, 50600,
  50600, 50601,
  50601, 50602,
  50602, 50603,
  50603, 50604,
  50604, 50605,
  50605, 50606,
  50606, 50607,
  50607, 50608,
  50608, 50609,
  50609, 50610,
  50610, 50611,
  50611, 50612,
  50612, 50613,
  50613, 50614,
  50614, 50615,
  50615, 50616,
  50616, 50617,
  50617, 50618,
  50618, 50619,
  50619, 50620,
  50620, 50621,
  50621, 50622,
  50622, 50623,
  50623, 50624,
  50624, 50625,
  50625, 50626,
  50626, 50627,
  50627, 50628,
  50628, 50629,
  50629, 50630,
  50630, 50631,
  50631, 50632,
  50632, 50633,
  50633, 50634,
  50634, 50635,
  50635, 50636,
  50636, 50637,
  50637, 50638,
  50638, 50639,
  50639, 50640,
  50640, 50641,
  50641, 50642,
  50642, 50643,
  50643, 50644,
  50644, 50645,
  50645, 50646,
  50646, 50647,
  50647, 50648,
  50648, 50649,
  50649, 50650,
  50650, 50651,
  50651, 50652,
  50652, 50653,
  50653, 50654,
  50654, 50655,
  50655, 50656,
  50656, 50657,
  50657, 50658,
  50658, 50659,
  50659, 50660,
  50660, 50661,
  50661, 50662,
  50662, 50663,
  50663, 50664,
  50664, 50665,
  50665, 50666,
  50666, 50667,
  50667, 50668,
  50668, 50669,
  50669, 50670,
  50670, 50671,
  50671, 50672,
  50672, 50673,
  50673, 50674,
  50674, 50675,
  50675, 50676,
  50676, 50677,
  50677, 50678,
  50678, 50679,
  50679, 50680,
  50680, 50681,
  50681, 50682,
  50682, 50683,
  50683, 50684,
  50684, 50685,
  50685, 50686,
  50686, 50687,
  50687, 50688,
  50688, 50689,
  50689, 50690,
  50690, 50691,
  50691, 50692,
  50692, 50693,
  50693, 50694,
  50694, 50695,
  50695, 50696,
  50696, 50697,
  50697, 50698,
  50698, 50699,
  50699, 50700,
  50700, 50701,
  50701, 50702,
  50702, 50703,
  50703, 50704,
  50704, 50705,
  50705, 50706,
  50706, 50707,
  50707, 50708,
  50708, 50709,
  50709, 50710,
  50710, 50711,
  50711, 50712,
  50712, 50713,
  50713, 50714,
  50714, 50715,
  50715, 50716,
  50716, 50717,
  50717, 50718,
  50718, 50719,
  50719, 50720,
  50720, 50721,
  50721, 50722,
  50722, 50723,
  50723, 50724,
  50724, 50725,
  50725, 50726,
  50726, 50727,
  50727, 50728,
  50728, 50729,
  50729, 50730,
  50730, 50731,
  50731, 50732,
  50732, 50733,
  50733, 50734,
  50734, 50735,
  50735, 50736,
  50736, 50737,
  50737, 50738,
  50738, 50739,
  50739, 50740,
  50740, 50741,
  50741, 50742,
  50742, 50743,
  50743, 50744,
  50744, 50745,
  50745, 50746,
  50746, 50747,
  50747, 50748,
  50748, 50749,
  50749, 50750,
  50750, 50751,
  50751, 50752,
  50752, 50753,
  50753, 50754,
  50754, 50755,
  50755, 50756,
  50756, 50757,
  50757, 50758,
  50758, 50759,
  50759, 50760,
  50760, 50761,
  50761, 50762,
  50762, 50763,
  50763, 50764,
  50764, 50765,
  50765, 50766,
  50766, 50767,
  50767, 50768,
  50768, 50769,
  50769, 50770,
  50770, 50771,
  50771, 50772,
  50772, 50773,
  50773, 50774,
  50774, 50775,
  50775, 50776,
  50776, 50777,
  50777, 50778,
  50778, 50779,
  50779, 50780,
  50780, 50781,
  50781, 50782,
  50782, 50783,
  50783, 50784,
  50784, 50785,
  50785, 50786,
  50786, 50787,
  50787, 50788,
  50788, 50789,
  50789, 50790,
  50790, 50791,
  50791, 50792,
  50792, 50793,
  50793, 50794,
  50794, 50795,
  50795, 50796,
  50796, 50797,
  50797, 50798,
  50798, 50799,
  50799, 50800,
  50800, 50801,
  50801, 50802,
  50802, 50803,
  50803, 50804,
  50804, 50805,
  50805, 50806,
  50806, 50807,
  50807, 50808,
  50808, 50809,
  50809, 50810,
  50810, 50811,
  50811, 50812,
  50812, 50813,
  50813, 50814,
  50814, 50815,
  50815, 50816,
  50816, 50817,
  50817, 50818,
  50818, 50819,
  50819, 50820,
  50820, 50821,
  50821, 50822,
  50822, 50823,
  50823, 50824,
  50824, 50825,
  50825, 50826,
  50826, 50827,
  50827, 50828,
  50828, 50829,
  50829, 50830,
  50830, 50831,
  50831, 50832,
  50832, 50833,
  50833, 50834,
  50834, 50835,
  50835, 50836,
  50836, 50837,
  50837, 50838,
  50838, 50839,
  50839, 50840,
  50840, 50841,
  50841, 50842,
  50842, 50843,
  50843, 50844,
  50844, 50845,
  50845, 50846,
  50846, 50847,
  50847, 50848,
  50848, 50849,
  50849, 50850,
  50850, 50851,
  50851, 50852,
  50852, 50853,
  50853, 50854,
  50854, 50855,
  50855, 50856,
  50856, 50857,
  50857, 50858,
  50858, 50859,
  50859, 50860,
  50860, 50861,
  50861, 50862,
  50862, 50863,
  50863, 50864,
  50864, 50865,
  50865, 50866,
  50866, 50867,
  50867, 50868,
  50868, 50869,
  50869, 50870,
  50870, 50871,
  50871, 50872,
  50872, 50873,
  50873, 50874,
  50874, 50875,
  50875, 50876,
  50876, 50877,
  50877, 50878,
  50878, 50879,
  50879, 50880,
  50880, 50881,
  50881, 50882,
  50882, 50883,
  50883, 50884,
  50884, 50885,
  50885, 50886,
  50886, 50887,
  50887, 50888,
  50888, 50889,
  50889, 50890,
  50890, 50891,
  50891, 50892,
  50892, 50893,
  50893, 50894,
  50894, 50895,
  50895, 50896,
  50896, 50897,
  50897, 50898,
  50898, 50899,
  50899, 50900,
  50900, 50901,
  50901, 50902,
  50902, 50903,
  50903, 50904,
  50904, 50905,
  50905, 50906,
  50906, 50907,
  50907, 50908,
  50908, 50909,
  50909, 50910,
  50910, 50911,
  50911, 50912,
  50912, 50913,
  50913, 50914,
  50914, 50915,
  50915, 50916,
  50916, 50917,
  50917, 50918,
  50918, 50919,
  50919, 50920,
  50920, 50921,
  50921, 50922,
  50922, 50923,
  50923, 50924,
  50924, 50925,
  50925, 50926,
  50926, 50927,
  50927, 50928,
  50928, 50929,
  50929, 50930,
  50930, 50931,
  50931, 50932,
  50932, 50933,
  50933, 50934,
  50934, 50935,
  50935, 50936,
  50936, 50937,
  50937, 50938,
  50938, 50939,
  50939, 50940,
  50940, 50941,
  50941, 50942,
  50942, 50943,
  50943, 50944,
  50944, 50945,
  50945, 50946,
  50946, 50947,
  50947, 50948,
  50948, 50949,
  50949, 50950,
  50950, 50951,
  50951, 50952,
  50952, 50953,
  50953, 50954,
  50954, 50955,
  50955, 50956,
  50956, 50957,
  50957, 50958,
  50958, 50959,
  50959, 50960,
  50960, 50961,
  50961, 50962,
  50962, 50963,
  50963, 50964,
  50964, 50965,
  50965, 50966,
  50966, 50967,
  50967, 50968,
  50968, 50969,
  50969, 50970,
  50970, 50971,
  50971, 50972,
  50972, 50973,
  50973, 50974,
  50974, 50975,
  50975, 50976,
  50976, 50977,
  50977, 50978,
  50978, 50979,
  50979, 50980,
  50980, 50981,
  50981, 50982,
  50982, 50983,
  50983, 50984,
  50984, 50985,
  50985, 50986,
  50986, 50987,
  50987, 50988,
  50988, 50989,
  50989, 50990,
  50990, 50991,
  50991, 50992,
  50992, 50993,
  50993, 50994,
  50994, 50995,
  50995, 50996,
  50996, 50997,
  50997, 50998,
  50998, 50999,
  50999, 51000,
  51000, 51001,
  51001, 51002,
  51002, 51003,
  51003, 51004,
  51004, 51005,
  51005, 51006,
  51006, 51007,
  51007, 51008,
  51008, 51009,
  51009, 51010,
  51010, 51011,
  51011, 51012,
  51012, 51013,
  51013, 51014,
  51014, 51015,
  51015, 51016,
  51016, 51017,
  51017, 51018,
  51018, 51019,
  51019, 51020,
  51020, 51021,
  51021, 51022,
  51022, 51023,
  51023, 51024,
  51024, 51025,
  51025, 51026,
  51026, 51027,
  51027, 51028,
  51028, 51029,
  51029, 51030,
  51030, 51031,
  51031, 51032,
  51032, 51033,
  51033, 51034,
  51034, 51035,
  51035, 51036,
  51036, 51037,
  51037, 51038,
  51038, 51039,
  51039, 51040,
  51040, 51041,
  51041, 51042,
  51042, 51043,
  51043, 51044,
  51044, 51045,
  51045, 51046,
  51046, 51047,
  51047, 51048,
  51048, 51049,
  51049, 51050,
  51050, 51051,
  51051, 51052,
  51052, 51053,
  51053, 51054,
  51054, 51055,
  51055, 51056,
  51056, 51057,
  51057, 51058,
  51058, 51059,
  51059, 51060,
  51060, 51061,
  51061, 51062,
  51062, 51063,
  51063, 51064,
  51064, 51065,
  51065, 51066,
  51066, 51067,
  51067, 51068,
  51068, 51069,
  51069, 51070,
  51070, 51071,
  51071, 51072,
  51072, 51073,
  51073, 51074,
  51074, 51075,
  51075, 51076,
  51076, 51077,
  51077, 51078,
  51078, 51079,
  51079, 51080,
  51080, 51081,
  51081, 51082,
  51082, 51083,
  51083, 51084,
  51084, 51085,
  51085, 51086,
  51086, 51087,
  51087, 51088,
  51088, 51089,
  51089, 51090,
  51090, 51091,
  51091, 51092,
  51092, 51093,
  51093, 51094,
  51094, 51095,
  51095, 51096,
  51096, 51097,
  51097, 51098,
  51098, 51099,
  51099, 51100,
  51100, 51101,
  51101, 51102,
  51102, 51103,
  51103, 51104,
  51104, 51105,
  51105, 51106,
  51106, 51107,
  51107, 51108,
  51108, 51109,
  51109, 51110,
  51110, 51111,
  51111, 51112,
  51112, 51113,
  51113, 51114,
  51114, 51115,
  51115, 51116,
  51116, 51117,
  51117, 51118,
  51118, 51119,
  51119, 51120,
  51120, 51121,
  51121, 51122,
  51122, 51123,
  51123, 51124,
  51124, 51125,
  51125, 51126,
  51126, 51127,
  51127, 51128,
  51128, 51129,
  51129, 51130,
  51130, 51131,
  51131, 51132,
  51132, 51133,
  51133, 51134,
  51134, 51135,
  51135, 51136,
  51136, 51137,
  51137, 51138,
  51138, 51139,
  51139, 51140,
  51140, 51141,
  51141, 51142,
  51142, 51143,
  51143, 51144,
  51144, 51145,
  51145, 51146,
  51146, 51147,
  51147, 51148,
  51148, 51149,
  51149, 51150,
  51150, 51151,
  51151, 51152,
  51152, 51153,
  51153, 51154,
  51154, 51155,
  51155, 51156,
  51156, 51157,
  51157, 51158,
  51158, 51159,
  51159, 51160,
  51160, 51161,
  51161, 51162,
  51162, 51163,
  51163, 51164,
  51164, 51165,
  51165, 51166,
  51166, 51167,
  51167, 51168,
  51168, 51169,
  51169, 51170,
  51170, 51171,
  51171, 51172,
  51172, 51173,
  51173, 51174,
  51174, 51175,
  51175, 51176,
  51176, 51177,
  51177, 51178,
  51178, 51179,
  51179, 51180,
  51180, 51181,
  51181, 51182,
  51182, 51183,
  51183, 51184,
  51184, 51185,
  51185, 51186,
  51186, 51187,
  51187, 51188,
  51188, 51189,
  51189, 51190,
  51190, 51191,
  51191, 51192,
  51192, 51193,
  51193, 51194,
  51194, 51195,
  51195, 51196,
  51196, 51197,
  51197, 51198,
  51198, 51199,
  51199, 51200,
  51200, 51201,
  51201, 51202,
  51202, 51203,
  51203, 51204,
  51204, 51205,
  51205, 51206,
  51206, 51207,
  51207, 51208,
  51208, 51209,
  51209, 51210,
  51210, 51211,
  51211, 51212,
  51212, 51213,
  51213, 51214,
  51214, 51215,
  51215, 51216,
  51216, 51217,
  51217, 51218,
  51218, 51219,
  51219, 51220,
  51220, 51221,
  51221, 51222,
  51222, 51223,
  51223, 51224,
  51224, 51225,
  51225, 51226,
  51226, 51227,
  51227, 51228,
  51228, 51229,
  51229, 51230,
  51230, 51231,
  51231, 51232,
  51232, 51233,
  51233, 51234,
  51234, 51235,
  51235, 51236,
  51236, 51237,
  51237, 51238,
  51238, 51239,
  51239, 51240,
  51240, 51241,
  51241, 51242,
  51242, 51243,
  51243, 51244,
  51244, 51245,
  51245, 51246,
  51246, 51247,
  51247, 51248,
  51248, 51249,
  51249, 51250,
  51250, 51251,
  51251, 51252,
  51252, 51253,
  51253, 51254,
  51254, 51255,
  51255, 51256,
  51256, 51257,
  51257, 51258,
  51258, 51259,
  51259, 51260,
  51260, 51261,
  51261, 51262,
  51262, 51263,
  51263, 51264,
  51264, 51265,
  51265, 51266,
  51266, 51267,
  51267, 51268,
  51268, 51269,
  51269, 51270,
  51270, 51271,
  51271, 51272,
  51272, 51273,
  51273, 51274,
  51274, 51275,
  51275, 51276,
  51276, 51277,
  51277, 51278,
  51278, 51279,
  51279, 51280,
  51280, 51281,
  51281, 51282,
  51282, 51283,
  51283, 51284,
  51284, 51285,
  51285, 51286,
  51286, 51287,
  51287, 51288,
  51288, 51289,
  51289, 51290,
  51290, 51291,
  51291, 51292,
  51292, 51293,
  51293, 51294,
  51294, 51295,
  51295, 51296,
  51296, 51297,
  51297, 51298,
  51298, 51299,
  51299, 51300,
  51300, 51301,
  51301, 51302,
  51302, 51303,
  51303, 51304,
  51304, 51305,
  51305, 51306,
  51306, 51307,
  51307, 51308,
  51308, 51309,
  51309, 51310,
  51310, 51311,
  51311, 51312,
  51312, 51313,
  51313, 51314,
  51314, 51315,
  51315, 51316,
  51316, 51317,
  51317, 51318,
  51318, 51319,
  51319, 51320,
  51320, 51321,
  51321, 51322,
  51322, 51323,
  51323, 51324,
  51324, 51325,
  51325, 51326,
  51326, 51327,
  51327, 51328,
  51328, 51329,
  51329, 51330,
  51330, 51331,
  51331, 51332,
  51332, 51333,
  51333, 51334,
  51334, 51335,
  51335, 51336,
  51336, 51337,
  51337, 51338,
  51338, 51339,
  51339, 51340,
  51340, 51341,
  51341, 51342,
  51342, 51343,
  51343, 51344,
  51344, 51345,
  51345, 51346,
  51346, 51347,
  51347, 51348,
  51348, 51349,
  51349, 51350,
  51350, 51351,
  51351, 51352,
  51352, 51353,
  51353, 51354,
  51354, 51355,
  51355, 51356,
  51356, 51357,
  51357, 51358,
  51358, 51359,
  51359, 51360,
  51360, 51361,
  51361, 51362,
  51362, 51363,
  51363, 51364,
  51364, 51365,
  51365, 51366,
  51366, 51367,
  51367, 51368,
  51368, 51369,
  51369, 51370,
  51370, 51371,
  51371, 51372,
  51372, 51373,
  51373, 51374,
  51374, 51375,
  51375, 51376,
  51376, 51377,
  51377, 51378,
  51378, 51379,
  51379, 51380,
  51380, 51381,
  51381, 51382,
  51382, 51383,
  51383, 51384,
  51384, 51385,
  51385, 51386,
  51386, 51387,
  51387, 51388,
  51388, 51389,
  51389, 51390,
  51390, 51391,
  51391, 51392,
  51392, 51393,
  51393, 51394,
  51394, 51395,
  51395, 51396,
  51396, 51397,
  51397, 51398,
  51398, 51399,
  51399, 51400,
  51400, 51401,
  51401, 51402,
  51402, 51403,
  51403, 51404,
  51404, 51405,
  51405, 51406,
  51406, 51407,
  51407, 51408,
  51408, 51409,
  51409, 51410,
  51410, 51411,
  51411, 51412,
  51412, 51413,
  51413, 51414,
  51414, 51415,
  51415, 51416,
  51416, 51417,
  51417, 51418,
  51418, 51419,
  51419, 51420,
  51420, 51421,
  51421, 51422,
  51422, 51423,
  51423, 51424,
  51424, 51425,
  51425, 51426,
  51426, 51427,
  51427, 51428,
  51428, 51429,
  51429, 51430,
  51430, 51431,
  51431, 51432,
  51432, 51433,
  51433, 51434,
  51434, 51435,
  51435, 51436,
  51436, 51437,
  51437, 51438,
  51438, 51439,
  51439, 51440,
  51440, 51441,
  51441, 51442,
  51442, 51443,
  51443, 51444,
  51444, 51445,
  51445, 51446,
  51446, 51447,
  51447, 51448,
  51448, 51449,
  51449, 51450,
  51450, 51451,
  51451, 51452,
  51452, 51453,
  51453, 51454,
  51454, 51455,
  51455, 51456,
  51456, 51457,
  51457, 51458,
  51458, 51459,
  51459, 51460,
  51460, 51461,
  51461, 51462,
  51462, 51463,
  51463, 51464,
  51464, 51465,
  51465, 51466,
  51466, 51467,
  51467, 51468,
  51468, 51469,
  51469, 51470,
  51470, 51471,
  51471, 51472,
  51472, 51473,
  51473, 51474,
  51474, 51475,
  51475, 51476,
  51476, 51477,
  51477, 51478,
  51478, 51479,
  51479, 51480,
  51480, 51481,
  51481, 51482,
  51482, 51483,
  51483, 51484,
  51484, 51485,
  51485, 51486,
  51486, 51487,
  51487, 51488,
  51488, 51489,
  51489, 51490,
  51490, 51491,
  51491, 51492,
  51492, 51493,
  51493, 51494,
  51494, 51495,
  51495, 51496,
  51496, 51497,
  51497, 51498,
  51498, 51499,
  51499, 51500,
  51500, 51501,
  51501, 51502,
  51502, 51503,
  51503, 51504,
  51504, 51505,
  51505, 51506,
  51506, 51507,
  51507, 51508,
  51508, 51509,
  51509, 51510,
  51510, 51511,
  51511, 51512,
  51512, 51513,
  51513, 51514,
  51514, 51515,
  51515, 51516,
  51516, 51517,
  51517, 51518,
  51518, 51519,
  51519, 51520,
  51520, 51521,
  51521, 51522,
  51522, 51523,
  51523, 51524,
  51524, 51525,
  51525, 51526,
  51526, 51527,
  51527, 51528,
  51528, 51529,
  51529, 51530,
  51530, 51531,
  51531, 51532,
  51532, 51533,
  51533, 51534,
  51534, 51535,
  51535, 51536,
  51536, 51537,
  51537, 51538,
  51538, 51539,
  51539, 51540,
  51540, 51541,
  51541, 51542,
  51542, 51543,
  51543, 51544,
  51544, 51545,
  51545, 51546,
  51546, 51547,
  51547, 51548,
  51548, 51549,
  51549, 51550,
  51550, 51551,
  51551, 51552,
  51552, 51553,
  51553, 51554,
  51554, 51555,
  51555, 51556,
  51556, 51557,
  51557, 51558,
  51558, 51559,
  51559, 51560,
  51560, 51561,
  51561, 51562,
  51562, 51563,
  51563, 51564,
  51564, 51565,
  51565, 51566,
  51566, 51567,
  51567, 51568,
  51568, 51569,
  51569, 51570,
  51570, 51571,
  51571, 51572,
  51572, 51573,
  51573, 51574,
  51574, 51575,
  51575, 51576,
  51576, 51577,
  51577, 51578,
  51578, 51579,
  51579, 51580,
  51580, 51581,
  51581, 51582,
  51582, 51583,
  51583, 51584,
  51584, 51585,
  51585, 51586,
  51586, 51587,
  51587, 51588,
  51588, 51589,
  51589, 51590,
  51590, 51591,
  51591, 51592,
  51592, 51593,
  51593, 51594,
  51594, 51595,
  51595, 51596,
  51596, 51597,
  51597, 51598,
  51598, 51599,
  51599, 51600,
  51600, 51601,
  51601, 51602,
  51602, 51603,
  51603, 51604,
  51604, 51605,
  51605, 51606,
  51606, 51607,
  51607, 51608,
  51608, 51609,
  51609, 51610,
  51610, 51611,
  51611, 51612,
  51612, 51613,
  51613, 51614,
  51614, 51615,
  51615, 51616,
  51616, 51617,
  51617, 51618,
  51618, 51619,
  51619, 51620,
  51620, 51621,
  51621, 51622,
  51622, 51623,
  51623, 51624,
  51624, 51625,
  51625, 51626,
  51626, 51627,
  51627, 51628,
  51628, 51629,
  51629, 51630,
  51630, 51631,
  51631, 51632,
  51632, 51633,
  51633, 51634,
  51634, 51635,
  51635, 51636,
  51636, 51637,
  51637, 51638,
  51638, 51639,
  51639, 51640,
  51640, 51641,
  51641, 51642,
  51642, 51643,
  51643, 51644,
  51644, 51645,
  51645, 51646,
  51646, 51647,
  51647, 51648,
  51648, 51649,
  51649, 51650,
  51650, 51651,
  51651, 51652,
  51652, 51653,
  51653, 51654,
  51654, 51655,
  51655, 51656,
  51656, 51657,
  51657, 51658,
  51658, 51659,
  51659, 51660,
  51660, 51661,
  51661, 51662,
  51662, 51663,
  51663, 51664,
  51664, 51665,
  51665, 51666,
  51666, 51667,
  51667, 51668,
  51668, 51669,
  51669, 51670,
  51670, 51671,
  51671, 51672,
  51672, 51673,
  51673, 51674,
  51674, 51675,
  51675, 51676,
  51676, 51677,
  51677, 51678,
  51678, 51679,
  51679, 51680,
  51680, 51681,
  51681, 51682,
  51682, 51683,
  51683, 51684,
  51684, 51685,
  51685, 51686,
  51686, 51687,
  51687, 51688,
  51688, 51689,
  51689, 51690,
  51690, 51691,
  51691, 51692,
  51692, 51693,
  51693, 51694,
  51694, 51695,
  51695, 51696,
  51696, 51697,
  51697, 51698,
  51698, 51699,
  51699, 51700,
  51700, 51701,
  51701, 51702,
  51702, 51703,
  51703, 51704,
  51704, 51705,
  51705, 51706,
  51706, 51707,
  51707, 51708,
  51708, 51709,
  51709, 51710,
  51710, 51711,
  51711, 51712,
  51712, 51713,
  51713, 51714,
  51714, 51715,
  51715, 51716,
  51716, 51717,
  51717, 51718,
  51718, 51719,
  51719, 51720,
  51720, 51721,
  51721, 51722,
  51722, 51723,
  51723, 51724,
  51724, 51725,
  51725, 51726,
  51726, 51727,
  51727, 51728,
  51728, 51729,
  51729, 51730,
  51730, 51731,
  51731, 51732,
  51732, 51733,
  51733, 51734,
  51734, 51735,
  51735, 51736,
  51736, 51737,
  51737, 51738,
  51738, 51739,
  51739, 51740,
  51740, 51741,
  51741, 51742,
  51742, 51743,
  51743, 51744,
  51744, 51745,
  51745, 51746,
  51746, 51747,
  51747, 51748,
  51748, 51749,
  51749, 51750,
  51750, 51751,
  51751, 51752,
  51752, 51753,
  51753, 51754,
  51754, 51755,
  51755, 51756,
  51756, 51757,
  51757, 51758,
  51758, 51759,
  51759, 51760,
  51760, 51761,
  51761, 51762,
  51762, 51763,
  51763, 51764,
  51764, 51765,
  51765, 51766,
  51766, 51767,
  51767, 51768,
  51768, 51769,
  51769, 51770,
  51770, 51771,
  51771, 51772,
  51772, 51773,
  51773, 51774,
  51774, 51775,
  51775, 51776,
  51776, 51777,
  51777, 51778,
  51778, 51779,
  51779, 51780,
  51780, 51781,
  51781, 51782,
  51782, 51783,
  51783, 51784,
  51784, 51785,
  51785, 51786,
  51786, 51787,
  51787, 51788,
  51788, 51789,
  51789, 51790,
  51790, 51791,
  51791, 51792,
  51792, 51793,
  51793, 51794,
  51794, 51795,
  51795, 51796,
  51796, 51797,
  51797, 51798,
  51798, 51799,
  51799, 51800,
  51800, 51801,
  51801, 51802,
  51802, 51803,
  51803, 51804,
  51804, 51805,
  51805, 51806,
  51806, 51807,
  51807, 51808,
  51808, 51809,
  51809, 51810,
  51810, 51811,
  51811, 51812,
  51812, 51813,
  51813, 51814,
  51814, 51815,
  51815, 51816,
  51816, 51817,
  51817, 51818,
  51818, 51819,
  51819, 51820,
  51820, 51821,
  51821, 51822,
  51822, 51823,
  51823, 51824,
  51824, 51825,
  51825, 51826,
  51826, 51827,
  51827, 51828,
  51828, 51829,
  51829, 51830,
  51830, 51831,
  51831, 51832,
  51832, 51833,
  51833, 51834,
  51834, 51835,
  51835, 51836,
  51836, 51837,
  51837, 51838,
  51838, 51839,
  51839, 51840,
  51840, 51841,
  51841, 51842,
  51842, 51843,
  51843, 51844,
  51844, 51845,
  51845, 51846,
  51846, 51847,
  51847, 51848,
  51848, 51849,
  51849, 51850,
  51850, 51851,
  51851, 51852,
  51852, 51853,
  51853, 51854,
  51854, 51855,
  51855, 51856,
  51856, 51857,
  51857, 51858,
  51858, 51859,
  51859, 51860,
  51860, 51861,
  51861, 51862,
  51862, 51863,
  51863, 51864,
  51864, 51865,
  51865, 51866,
  51866, 51867,
  51867, 51868,
  51868, 51869,
  51869, 51870,
  51870, 51871,
  51871, 51872,
  51872, 51873,
  51873, 51874,
  51874, 51875,
  51875, 51876,
  51876, 51877,
  51877, 51878,
  51878, 51879,
  51879, 51880,
  51880, 51881,
  51881, 51882,
  51882, 51883,
  51883, 51884,
  51884, 51885,
  51885, 51886,
  51886, 51887,
  51887, 51888,
  51888, 51889,
  51889, 51890,
  51890, 51891,
  51891, 51892,
  51892, 51893,
  51893, 51894,
  51894, 51895,
  51895, 51896,
  51896, 51897,
  51897, 51898,
  51898, 51899,
  51899, 51900,
  51900, 51901,
  51901, 51902,
  51902, 51903,
  51903, 51904,
  51904, 51905,
  51905, 51906,
  51906, 51907,
  51907, 51908,
  51908, 51909,
  51909, 51910,
  51910, 51911,
  51911, 51912,
  51912, 51913,
  51913, 51914,
  51914, 51915,
  51915, 51916,
  51916, 51917,
  51917, 51918,
  51918, 51919,
  51919, 51920,
  51920, 51921,
  51921, 51922,
  51922, 51923,
  51923, 51924,
  51924, 51925,
  51925, 51926,
  51926, 51927,
  51927, 51928,
  51928, 51929,
  51929, 51930,
  51930, 51931,
  51931, 51932,
  51932, 51933,
  51933, 51934,
  51934, 51935,
  51935, 51936,
  51936, 51937,
  51937, 51938,
  51938, 51939,
  51939, 51940,
  51940, 51941,
  51941, 51942,
  51942, 51943,
  51943, 51944,
  51944, 51945,
  51945, 51946,
  51946, 51947,
  51947, 51948,
  51948, 51949,
  51949, 51950,
  51950, 51951,
  51951, 51952,
  51952, 51953,
  51953, 51954,
  51954, 51955,
  51955, 51956,
  51956, 51957,
  51957, 51958,
  51958, 51959,
  51959, 51960,
  51960, 51961,
  51961, 51962,
  51962, 51963,
  51963, 51964,
  51964, 51965,
  51965, 51966,
  51966, 51967,
  51967, 51968,
  51968, 51969,
  51969, 51970,
  51970, 51971,
  51971, 51972,
  51972, 51973,
  51973, 51974,
  51974, 51975,
  51975, 51976,
  51976, 51977,
  51977, 51978,
  51978, 51979,
  51979, 51980,
  51980, 51981,
  51981, 51982,
  51982, 51983,
  51983, 51984,
  51984, 51985,
  51985, 51986,
  51986, 51987,
  51987, 51988,
  51988, 51989,
  51989, 51990,
  51990, 51991,
  51991, 51992,
  51992, 51993,
  51993, 51994,
  51994, 51995,
  51995, 51996,
  51996, 51997,
  51997, 51998,
  51998, 51999,
  51999, 52000,
  52000, 52001,
  52001, 52002,
  52002, 52003,
  52003, 52004,
  52004, 52005,
  52005, 52006,
  52006, 52007,
  52007, 52008,
  52008, 52009,
  52009, 52010,
  52010, 52011,
  52011, 52012,
  52012, 52013,
  52013, 52014,
  52014, 52015,
  52015, 52016,
  52016, 52017,
  52017, 52018,
  52018, 52019,
  52019, 52020,
  52020, 52021,
  52021, 52022,
  52022, 52023,
  52023, 52024,
  52024, 52025,
  52025, 52026,
  52026, 52027,
  52027, 52028,
  52028, 52029,
  52029, 52030,
  52030, 52031,
  52031, 52032,
  52032, 52033,
  52033, 52034,
  52034, 52035,
  52035, 52036,
  52036, 52037,
  52037, 52038,
  52038, 52039,
  52039, 52040,
  52040, 52041,
  52041, 52042,
  52042, 52043,
  52043, 52044,
  52044, 52045,
  52045, 52046,
  52046, 52047,
  52047, 52048,
  52048, 52049,
  52049, 52050,
  52050, 52051,
  52051, 52052,
  52052, 52053,
  52053, 52054,
  52054, 52055,
  52055, 52056,
  52056, 52057,
  52057, 52058,
  52058, 52059,
  52059, 52060,
  52060, 52061,
  52061, 52062,
  52062, 52063,
  52063, 52064,
  52064, 52065,
  52065, 52066,
  52066, 52067,
  52067, 52068,
  52068, 52069,
  52069, 52070,
  52070, 52071,
  52071, 52072,
  52072, 52073,
  52073, 52074,
  52074, 52075,
  52075, 52076,
  52076, 52077,
  52077, 52078,
  52078, 52079,
  52079, 52080,
  52080, 52081,
  52081, 52082,
  52082, 52083,
  52083, 52084,
  52084, 52085,
  52085, 52086,
  52086, 52087,
  52087, 52088,
  52088, 52089,
  52089, 52090,
  52090, 52091,
  52091, 52092,
  52092, 52093,
  52093, 52094,
  52094, 52095,
  52095, 52096,
  52096, 52097,
  52097, 52098,
  52098, 52099,
  52099, 52100,
  52100, 52101,
  52101, 52102,
  52102, 52103,
  52103, 52104,
  52104, 52105,
  52105, 52106,
  52106, 52107,
  52107, 52108,
  52108, 52109,
  52109, 52110,
  52110, 52111,
  52111, 52112,
  52112, 52113,
  52113, 52114,
  52114, 52115,
  52115, 52116,
  52116, 52117,
  52117, 52118,
  52118, 52119,
  52119, 52120,
  52120, 52121,
  52121, 52122,
  52122, 52123,
  52123, 52124,
  52124, 52125,
  52125, 52126,
  52126, 52127,
  52127, 52128,
  52128, 52129,
  52129, 52130,
  52130, 52131,
  52131, 52132,
  52132, 52133,
  52133, 52134,
  52134, 52135,
  52135, 52136,
  52136, 52137,
  52137, 52138,
  52138, 52139,
  52139, 52140,
  52140, 52141,
  52141, 52142,
  52142, 52143,
  52143, 52144,
  52144, 52145,
  52145, 52146,
  52146, 52147,
  52147, 52148,
  52148, 52149,
  52149, 52150,
  52150, 52151,
  52151, 52152,
  52152, 52153,
  52153, 52154,
  52154, 52155,
  52155, 52156,
  52156, 52157,
  52157, 52158,
  52158, 52159,
  52159, 52160,
  52160, 52161,
  52161, 52162,
  52162, 52163,
  52163, 52164,
  52164, 52165,
  52165, 52166,
  52166, 52167,
  52167, 52168,
  52168, 52169,
  52169, 52170,
  52170, 52171,
  52171, 52172,
  52172, 52173,
  52173, 52174,
  52174, 52175,
  52175, 52176,
  52176, 52177,
  52177, 52178,
  52178, 52179,
  52179, 52180,
  52180, 52181,
  52181, 52182,
  52182, 52183,
  52183, 52184,
  52184, 52185,
  52185, 52186,
  52186, 52187,
  52187, 52188,
  52188, 52189,
  52189, 52190,
  52190, 52191,
  52191, 52192,
  52192, 52193,
  52193, 52194,
  52194, 52195,
  52195, 52196,
  52196, 52197,
  52197, 52198,
  52198, 52199,
  52199, 52200,
  52200, 52201,
  52201, 52202,
  52202, 52203,
  52203, 52204,
  52204, 52205,
  52205, 52206,
  52206, 52207,
  52207, 52208,
  52208, 52209,
  52209, 52210,
  52210, 52211,
  52211, 52212,
  52212, 52213,
  52213, 52214,
  52214, 52215,
  52215, 52216,
  52216, 52217,
  52217, 52218,
  52218, 52219,
  52219, 52220,
  52220, 52221,
  52221, 52222,
  52222, 52223,
  52223, 52224,
  52224, 52225,
  52225, 52226,
  52226, 52227,
  52227, 52228,
  52228, 52229,
  52229, 52230,
  52230, 52231,
  52231, 52232,
  52232, 52233,
  52233, 52234,
  52234, 52235,
  52235, 52236,
  52236, 52237,
  52237, 52238,
  52238, 52239,
  52239, 52240,
  52240, 52241,
  52241, 52242,
  52242, 52243,
  52243, 52244,
  52244, 52245,
  52245, 52246,
  52246, 52247,
  52247, 52248,
  52248, 52249,
  52249, 52250,
  52250, 52251,
  52251, 52252,
  52252, 52253,
  52253, 52254,
  52254, 52255,
  52255, 52256,
  52256, 52257,
  52257, 52258,
  52258, 52259,
  52259, 52260,
  52260, 52261,
  52261, 52262,
  52262, 52263,
  52263, 52264,
  52264, 52265,
  52265, 52266,
  52266, 52267,
  52267, 52268,
  52268, 52269,
  52269, 52270,
  52270, 52271,
  52271, 52272,
  52272, 52273,
  52273, 52274,
  52274, 52275,
  52275, 52276,
  52276, 52277,
  52277, 52278,
  52278, 52279,
  52279, 52280,
  52280, 52281,
  52281, 52282,
  52282, 52283,
  52283, 52284,
  52284, 52285,
  52285, 52286,
  52286, 52287,
  52287, 52288,
  52288, 52289,
  52289, 52290,
  52290, 52291,
  52291, 52292,
  52292, 52293,
  52293, 52294,
  52294, 52295,
  52295, 52296,
  52296, 52297,
  52297, 52298,
  52298, 52299,
  52299, 52300,
  52300, 52301,
  52301, 52302,
  52302, 52303,
  52303, 52304,
  52304, 52305,
  52305, 52306,
  52306, 52307,
  52307, 52308,
  52308, 52309,
  52309, 52310,
  52310, 52311,
  52311, 52312,
  52312, 52313,
  52313, 52314,
  52314, 52315,
  52315, 52316,
  52316, 52317,
  52317, 52318,
  52318, 52319,
  52319, 52320,
  52320, 52321,
  52321, 52322,
  52322, 52323,
  52323, 52324,
  52324, 52325,
  52325, 52326,
  52326, 52327,
  52327, 52328,
  52328, 52329,
  52329, 52330,
  52330, 52331,
  52331, 52332,
  52332, 52333,
  52333, 52334,
  52334, 52335,
  52335, 52336,
  52336, 52337,
  52337, 52338,
  52338, 52339,
  52339, 52340,
  52340, 52341,
  52341, 52342,
  52342, 52343,
  52343, 52344,
  52344, 52345,
  52345, 52346,
  52346, 52347,
  52347, 52348,
  52348, 52349,
  52349, 52350,
  52350, 52351,
  52351, 52352,
  52352, 52353,
  52353, 52354,
  52354, 52355,
  52355, 52356,
  52356, 52357,
  52357, 52358,
  52358, 52359,
  52359, 52360,
  52360, 52361,
  52361, 52362,
  52362, 52363,
  52363, 52364,
  52364, 52365,
  52365, 52366,
  52366, 52367,
  52367, 52368,
  52368, 52369,
  52369, 52370,
  52370, 52371,
  52371, 52372,
  52372, 52373,
  52373, 52374,
  52374, 52375,
  52375, 52376,
  52376, 52377,
  52377, 52378,
  52378, 52379,
  52379, 52380,
  52380, 52381,
  52381, 52382,
  52382, 52383,
  52383, 52384,
  52384, 52385,
  52385, 52386,
  52386, 52387,
  52387, 52388,
  52388, 52389,
  52389, 52390,
  52390, 52391,
  52391, 52392,
  52392, 52393,
  52393, 52394,
  52394, 52395,
  52395, 52396,
  52396, 52397,
  52397, 52398,
  52398, 52399,
  52399, 52400,
  52400, 52401,
  52401, 52402,
  52402, 52403,
  52403, 52404,
  52404, 52405,
  52405, 52406,
  52406, 52407,
  52407, 52408,
  52408, 52409,
  52409, 52410,
  52410, 52411,
  52411, 52412,
  52412, 52413,
  52413, 52414,
  52414, 52415,
  52415, 52416,
  52416, 52417,
  52417, 52418,
  52418, 52419,
  52419, 52420,
  52420, 52421,
  52421, 52422,
  52422, 52423,
  52423, 52424,
  52424, 52425,
  52425, 52426,
  52426, 52427,
  52427, 52428,
  52428, 52429,
  52429, 52430,
  52430, 52431,
  52431, 52432,
  52432, 52433,
  52433, 52434,
  52434, 52435,
  52435, 52436,
  52436, 52437,
  52437, 52438,
  52438, 52439,
  52439, 52440,
  52440, 52441,
  52441, 52442,
  52442, 52443,
  52443, 52444,
  52444, 52445,
  52445, 52446,
  52446, 52447,
  52447, 52448,
  52448, 52449,
  52449, 52450,
  52450, 52451,
  52451, 52452,
  52452, 52453,
  52453, 52454,
  52454, 52455,
  52455, 52456,
  52456, 52457,
  52457, 52458,
  52458, 52459,
  52459, 52460,
  52460, 52461,
  52461, 52462,
  52462, 52463,
  52463, 52464,
  52464, 52465,
  52465, 52466,
  52466, 52467,
  52467, 52468,
  52468, 52469,
  52469, 52470,
  52470, 52471,
  52471, 52472,
  52472, 52473,
  52473, 52474,
  52474, 52475,
  52475, 52476,
  52476, 52477,
  52477, 52478,
  52478, 52479,
  52479, 52480,
  52480, 52481,
  52481, 52482,
  52482, 52483,
  52483, 52484,
  52484, 52485,
  52485, 52486,
  52486, 52487,
  52487, 52488,
  52488, 52489,
  52489, 52490,
  52490, 52491,
  52491, 52492,
  52492, 52493,
  52493, 52494,
  52494, 52495,
  52495, 52496,
  52496, 52497,
  52497, 52498,
  52498, 52499,
  52499, 52500,
  52500, 52501,
  52501, 52502,
  52502, 52503,
  52503, 52504,
  52504, 52505,
  52505, 52506,
  52506, 52507,
  52507, 52508,
  52508, 52509,
  52509, 52510,
  52510, 52511,
  52511, 52512,
  52512, 52513,
  52513, 52514,
  52514, 52515,
  52515, 52516,
  52516, 52517,
  52517, 52518,
  52518, 52519,
  52519, 52520,
  52520, 52521,
  52521, 52522,
  52522, 52523,
  52523, 52524,
  52524, 52525,
  52525, 52526,
  52526, 52527,
  52527, 52528,
  52528, 52529,
  52529, 52530,
  52530, 52531,
  52531, 52532,
  52532, 52533,
  52533, 52534,
  52534, 52535,
  52535, 52536,
  52536, 52537,
  52537, 52538,
  52538, 52539,
  52539, 52540,
  52540, 52541,
  52541, 52542,
  52542, 52543,
  52543, 52544,
  52544, 52545,
  52545, 52546,
  52546, 52547,
  52547, 52548,
  52548, 52549,
  52549, 52550,
  52550, 52551,
  52551, 52552,
  52552, 52553,
  52553, 52554,
  52554, 52555,
  52555, 52556,
  52556, 52557,
  52557, 52558,
  52558, 52559,
  52559, 52560 ;
}
